module GLYPH_ROM2(piece, addr, row, value);
input [15:0]piece;
input [5:0] row;
input [5:0] addr;
output reg [0:39] value;

reg sqcolor;
//peice numbers
parameter  square = 3'b000 ,  pawn =3'b001 , rook = 3'b010 , horse = 3'b011, bishop = 3'b100, queen = 3'b101, king = 3'b110; 
//square color selection
always@(addr)begin
	if(addr <= 7 || (addr>= 16 && addr <= 23)//for the checkered pattern of the board 
	|| (addr>= 32 && addr <= 39) || (addr>= 48 && addr <= 55))begin
		if(addr % 2)
			sqcolor <= 0;//black square 
		else
			sqcolor <= 1;//white square
	end
	else begin
		if(addr % 2)
			sqcolor <= 1;//white square 
		else
			sqcolor <= 0;//black square 
	end


end


always@(*) begin

	//glyph selection
	case(piece[2:0])
		square: begin
			if(sqcolor)begin
				 case(row)//white square 
					0: value =  40'b1111111111111111111111111111111111111111;
					1: value =  40'b1111111111111111111111111111111111111111;
					2: value =  40'b1111111111111111111111111111111111111111;
					3: value =  40'b1111111111111111111111111111111111111111;
					4: value =  40'b1111111111111111111111111111111111111111;
					5: value =  40'b1111111111111111111111111111111111111111;
					6: value =  40'b1111111111111111111111111111111111111111;
					7: value =  40'b1111111111111111111111111111111111111111;
					8: value =  40'b1111111111111111111111111111111111111111;
					9: value =  40'b1111111111111111111111111111111111111111;
					10: value=  40'b1111111111111111111111111111111111111111;
					11: value = 40'b1111111111111111111111111111111111111111;
					12: value = 40'b1111111111111111111111111111111111111111;
					13: value = 40'b1111111111111111111111111111111111111111;
					14: value = 40'b1111111111111111111111111111111111111111;
					15: value = 40'b1111111111111111111111111111111111111111;
					16: value = 40'b1111111111111111111111111111111111111111;
					17: value = 40'b1111111111111111111111111111111111111111;
					18: value = 40'b1111111111111111111111111111111111111111;
					19: value = 40'b1111111111111111111111111111111111111111;
					20: value = 40'b1111111111111111111111111111111111111111;
					21: value = 40'b1111111111111111111111111111111111111111;
					22: value = 40'b1111111111111111111111111111111111111111;
					23: value = 40'b1111111111111111111111111111111111111111;
					24: value = 40'b1111111111111111111111111111111111111111;
					25: value = 40'b1111111111111111111111111111111111111111;
					26: value = 40'b1111111111111111111111111111111111111111;
					27: value = 40'b1111111111111111111111111111111111111111;
					28: value = 40'b1111111111111111111111111111111111111111;
					29: value = 40'b1111111111111111111111111111111111111111;
					30: value = 40'b1111111111111111111111111111111111111111;
					31: value = 40'b1111111111111111111111111111111111111111;
					32: value = 40'b1111111111111111111111111111111111111111;
					33: value = 40'b1111111111111111111111111111111111111111;
					34: value = 40'b1111111111111111111111111111111111111111;
					35: value = 40'b1111111111111111111111111111111111111111;
					36: value = 40'b1111111111111111111111111111111111111111;
					37: value = 40'b1111111111111111111111111111111111111111;
					38: value = 40'b1111111111111111111111111111111111111111;
					39: value = 40'b1111111111111111111111111111111111111111;
					default: value = 40'd0;
				endcase 
					
			end
			else begin
				 case(row) //black square
					0: value =  40'b0000000000000000000000000000000000000000;
					1: value =  40'b0000000000000000000000000000000000000000;
					2: value =  40'b0000000000000000000000000000000000000000;
					3: value =  40'b0000000000000000000000000000000000000000;
					4: value =  40'b0000000000000000000000000000000000000000;
					5: value =  40'b0000000000000000000000000000000000000000;
					6: value =  40'b0000000000000000000000000000000000000000;
					7: value =  40'b0000000000000000000000000000000000000000;
					8: value =  40'b0000000000000000000000000000000000000000;
					9: value =  40'b0000000000000000000000000000000000000000;
					10: value=  40'b0000000000000000000000000000000000000000;
					11: value = 40'b0000000000000000000000000000000000000000;
					12: value = 40'b0000000000000000000000000000000000000000;
					13: value = 40'b0000000000000000000000000000000000000000;
					14: value = 40'b0000000000000000000000000000000000000000;
					15: value = 40'b0000000000000000000000000000000000000000;
					16: value = 40'b0000000000000000000000000000000000000000;
					17: value = 40'b0000000000000000000000000000000000000000;
					18: value = 40'b0000000000000000000000000000000000000000;
					19: value = 40'b0000000000000000000000000000000000000000;
					20: value = 40'b0000000000000000000000000000000000000000;
					21: value = 40'b0000000000000000000000000000000000000000;
					22: value = 40'b0000000000000000000000000000000000000000;
					23: value = 40'b0000000000000000000000000000000000000000;
					24: value = 40'b0000000000000000000000000000000000000000;
					25: value = 40'b0000000000000000000000000000000000000000;
					26: value = 40'b0000000000000000000000000000000000000000;
					27: value = 40'b0000000000000000000000000000000000000000;
					28: value = 40'b0000000000000000000000000000000000000000;
					29: value = 40'b0000000000000000000000000000000000000000;
					30: value = 40'b0000000000000000000000000000000000000000;
					31: value = 40'b0000000000000000000000000000000000000000;
					32: value = 40'b0000000000000000000000000000000000000000;
					33: value = 40'b0000000000000000000000000000000000000000;
					34: value = 40'b0000000000000000000000000000000000000000;
					35: value = 40'b0000000000000000000000000000000000000000;
					36: value = 40'b0000000000000000000000000000000000000000;
					37: value = 40'b0000000000000000000000000000000000000000;
					38: value = 40'b0000000000000000000000000000000000000000;
					39: value = 40'b0000000000000000000000000000000000000000;
					default: value = 40'd0;
				endcase 
			
			end
		
		end
		
		pawn:begin
			if(piece > 7)begin // if piece is white or black
				if(sqcolor)begin
					case(row)//white square white pawn
			0: value =  40'b1111111111111111111111111111111111111111;
			1: value =  40'b1111111111111111111111111111111111111111;
			2: value =  40'b1111111111111111111111111111111111111111;
			3: value =  40'b1111111111111111111111111111111111111111;
			4: value =  40'b1111111111111111100000011111111111111111;
			5: value =  40'b1111111111111111011111101111111111111111;
			6: value =  40'b1111111111111110111111110111111111111111;
			7: value =  40'b1111111111111101111111111011111111111111;
			8: value =  40'b1111111111111101111111111011111111111111;
			9: value =  40'b1111111111111101111111111011111111111111;
			10: value=  40'b1111111111111110111111110111111111111111;
			11: value = 40'b1111111111111111011111101111111111111111;
			12: value = 40'b1111111111111110111111110111111111111111;
			13: value = 40'b1111111111111101111111111011111111111111;
			14: value = 40'b1111111111111011111111111101111111111111;
			15: value = 40'b1111111111110111111111111110111111111111;
			16: value = 40'b1111111111110111111111111110111111111111;
			17: value = 40'b1111111111110111111111111110111111111111;
			18: value = 40'b1111111111110111111111111110111111111111;
			19: value = 40'b1111111111111011111111111101111111111111;
			20: value = 40'b1111111111111101111111111011111111111111;
			21: value = 40'b1111111111111110111111110111111111111111;
			22: value = 40'b1111111111111111011111101111111111111111;
			23: value = 40'b1111111111111110111111110111111111111111;
			24: value = 40'b1111111111111101111111111011111111111111;
			25: value = 40'b1111111111111011111111111101111111111111;
			26: value = 40'b1111111111110111111111111110111111111111;
			27: value = 40'b1111111111101111111111111111011111111111;
			28: value = 40'b1111111111011111111111111111101111111111;
			29: value = 40'b1111111110111111111111111111110111111111;
			30: value = 40'b1111111101111111111111111111111011111111;
			31: value = 40'b1111111011111111111111111111111101111111;
			32: value = 40'b1111110111111111111111111111111110111111;
			33: value = 40'b1111101111111111111111111111111111011111;
			34: value = 40'b1111101111111111111111111111111111011111;
			35: value = 40'b1111100000000000000000000000000000011111;
			36: value = 40'b1111111111111111111111111111111111111111;
			37: value = 40'b1111111111111111111111111111111111111111;
			38: value = 40'b1111111111111111111111111111111111111111;
			39: value = 40'b1111111111111111111111111111111111111111;
			default: value = 40'd0;
		endcase 

				
				end
				else begin
					case(row) //black square white pawn
			0: value =  40'b0000000000000000000000000000000000000000;
			1: value =  40'b0000000000000000000000000000000000000000;
			2: value =  40'b0000000000000000000000000000000000000000;
			3: value =  40'b0000000000000000000000000000000000000000;
			4: value =  40'b0000000000000000000000000000000000000000;
			5: value =  40'b0000000000000000011111100000000000000000;
			6: value =  40'b0000000000000000111111110000000000000000;
			7: value =  40'b0000000000000001111111111000000000000000;
			8: value =  40'b0000000000000001111111111000000000000000;
			9: value =  40'b0000000000000001111111111000000000000000;
			10: value=  40'b0000000000000000111111110000000000000000;
			11: value = 40'b0000000000000000011111100000000000000000;
			12: value = 40'b0000000000000000111111110000000000000000;
			13: value = 40'b0000000000000001111111111000000000000000;
			14: value = 40'b0000000000000011111111111100000000000000;
			15: value = 40'b0000000000000111111111111110000000000000;
			16: value = 40'b0000000000000111111111111110000000000000;
			17: value = 40'b0000000000000111111111111110000000000000;
			18: value = 40'b0000000000000111111111111110000000000000;
			19: value = 40'b0000000000000011111111111100000000000000;
			20: value = 40'b0000000000000001111111111000000000000000;
			21: value = 40'b0000000000000000111111110000000000000000;
			22: value = 40'b0000000000000000011111100000000000000000;
			23: value = 40'b0000000000000000111111110000000000000000;
			24: value = 40'b0000000000000001111111111000000000000000;
			25: value = 40'b0000000000000011111111111100000000000000;
			26: value = 40'b0000000000000111111111111110000000000000;
			27: value = 40'b0000000000001111111111111111000000000000;
			28: value = 40'b0000000000011111111111111111100000000000;
			29: value = 40'b0000000000111111111111111111110000000000;
			30: value = 40'b0000000001111111111111111111111000000000;
			31: value = 40'b0000000011111111111111111111111100000000;
			32: value = 40'b0000000111111111111111111111111110000000;
			33: value = 40'b0000001111111111111111111111111111000000;
			34: value = 40'b0000001111111111111111111111111111000000;
			35: value = 40'b0000000000000000000000000000000000000000;
			36: value = 40'b0000000000000000000000000000000000000000;
			37: value = 40'b0000000000000000000000000000000000000000;
			38: value = 40'b0000000000000000000000000000000000000000;
			39: value = 40'b0000000000000000000000000000000000000000;
			default: value = 40'd0;
		endcase 

				end
			end
			else begin
				if(sqcolor)begin
					case(row)//white square black pawn
			0: value =  40'b1111111111111111111111111111111111111111;
			1: value =  40'b1111111111111111111111111111111111111111;
			2: value =  40'b1111111111111111111111111111111111111111;
			3: value =  40'b1111111111111111111111111111111111111111;
			4: value =  40'b1111111111111111111111111111111111111111;
			5: value =  40'b1111111111111111100000011111111111111111;
			6: value =  40'b1111111111111111000000001111111111111111;
			7: value =  40'b1111111111111110000000000111111111111111;
			8: value =  40'b1111111111111110000000000111111111111111;
			9: value =  40'b1111111111111110000000000111111111111111;
			10: value=  40'b1111111111111111000000001111111111111111;
			11: value = 40'b1111111111111111100000011111111111111111;
			12: value = 40'b1111111111111111000000001111111111111111;
			13: value = 40'b1111111111111110000000000111111111111111;
			14: value = 40'b1111111111111100000000000011111111111111;
			15: value = 40'b1111111111111000000000000001111111111111;
			16: value = 40'b1111111111111000000000000001111111111111;
			17: value = 40'b1111111111111000000000000001111111111111;
			18: value = 40'b1111111111111000000000000001111111111111;
			19: value = 40'b1111111111111100000000000011111111111111;
			20: value = 40'b1111111111111110000000000111111111111111;
			21: value = 40'b1111111111111111000000001111111111111111;
			22: value = 40'b1111111111111111100000011111111111111111;
			23: value = 40'b1111111111111111000000001111111111111111;
			24: value = 40'b1111111111111110000000000111111111111111;
			25: value = 40'b1111111111111100000000000011111111111111;
			26: value = 40'b1111111111111000000000000001111111111111;
			27: value = 40'b1111111111110000000000000000111111111111;
			28: value = 40'b1111111111100000000000000000011111111111;
			29: value = 40'b1111111111000000000000000000001111111111;
			30: value = 40'b1111111110000000000000000000000111111111;
			31: value = 40'b1111111100000000000000000000000011111111;
			32: value = 40'b1111111000000000000000000000000001111111;
			33: value = 40'b1111110000000000000000000000000000111111;
			34: value = 40'b1111110000000000000000000000000000111111;
			35: value = 40'b1111111111111111111111111111111111111111;
			36: value = 40'b1111111111111111111111111111111111111111;
			37: value = 40'b1111111111111111111111111111111111111111;
			38: value = 40'b1111111111111111111111111111111111111111;
			39: value = 40'b1111111111111111111111111111111111111111;
			default: value = 40'd0;
		endcase 
				
				end
				else begin
					case(row) //black square black pawn
			0: value =  40'b0000000000000000000000000000000000000000;
			1: value =  40'b0000000000000000000000000000000000000000;
			2: value =  40'b0000000000000000000000000000000000000000;
			3: value =  40'b0000000000000000000000000000000000000000;
			4: value =  40'b0000000000000000011111100000000000000000;
			5: value =  40'b0000000000000000100000010000000000000000;
			6: value =  40'b0000000000000001000000001000000000000000;
			7: value =  40'b0000000000000010000000000100000000000000;
			8: value =  40'b0000000000000010000000000100000000000000;
			9: value =  40'b0000000000000010000000000100000000000000;
			10: value=  40'b0000000000000001000000001000000000000000;
			11: value = 40'b0000000000000000100000010000000000000000;
			12: value = 40'b0000000000000001000000001000000000000000;
			13: value = 40'b0000000000000010000000000100000000000000;
			14: value = 40'b0000000000000100000000000010000000000000;
			15: value = 40'b0000000000001000000000000001000000000000;
			16: value = 40'b0000000000001000000000000001000000000000;
			17: value = 40'b0000000000001000000000000001000000000000;
			18: value = 40'b0000000000001000000000000001000000000000;
			19: value = 40'b0000000000000100000000000010000000000000;
			20: value = 40'b0000000000000010000000000100000000000000;
			21: value = 40'b0000000000000001000000001000000000000000;
			22: value = 40'b0000000000000000100000010000000000000000;
			23: value = 40'b0000000000000001000000001000000000000000;
			24: value = 40'b0000000000000010000000000100000000000000;
			25: value = 40'b0000000000000100000000000010000000000000;
			26: value = 40'b0000000000001000000000000001000000000000;
			27: value = 40'b0000000000010000000000000000100000000000;
			28: value = 40'b0000000000100000000000000000010000000000;
			29: value = 40'b0000000001000000000000000000001000000000;
			30: value = 40'b0000000010000000000000000000000100000000;
			31: value = 40'b0000000100000000000000000000000010000000;
			32: value = 40'b0000001000000000000000000000000001000000;
			33: value = 40'b0000010000000000000000000000000000100000;
			34: value = 40'b0000010000000000000000000000000000100000;
			35: value = 40'b0000011111111111111111111111111111100000;
			36: value = 40'b0000000000000000000000000000000000000000;
			37: value = 40'b0000000000000000000000000000000000000000;
			38: value = 40'b0000000000000000000000000000000000000000;
			39: value = 40'b0000000000000000000000000000000000000000;
			default: value = 40'd0;
		endcase 

				end
			end
		end
		
		rook:begin
			if(piece > 7)begin // if piece is white or black
				if(sqcolor)begin
						case(row)//white square white rook
			0: value =  40'b1111111111111111111111111111111111111111;
			1: value =  40'b1111111111111111111111111111111111111111;
			2: value =  40'b1111111111111111111111111111111111111111;
			3: value =  40'b1111111111111111111111111111111111111111;
			4: value =  40'b1111100000000010000000000100000000011111;
			5: value =  40'b1111101111111010111111110101111111011111;
			6: value =  40'b1111101111111010111111110101111111011111;
			7: value =  40'b1111101111111010111111110101111111011111;
			8: value =  40'b1111101111111000111111110001111111011111;
			9: value=   40'b1111101111111111111111111111111111011111;
			10: value = 40'b1111101111111111111111111111111111011111;
			11: value = 40'b1111101111111111111111111111111111011111;
			12: value = 40'b1111101111111111111111111111111111011111;
			13: value = 40'b1111101111111111111111111111111111011111;
			14: value = 40'b1111101111111111111111111111111111011111;
			15: value = 40'b1111101111111111111111111111111111011111;
			16: value = 40'b1111100000001111111111111111000000011111;
			17: value = 40'b1111111111101111111111111111011111111111;
			18: value = 40'b1111111111101111111111111111011111111111;
			19: value = 40'b1111111000001111111111111111000001111111;
			20: value = 40'b1111111011111111111111111111111101111111;
			21: value = 40'b1111111011111111111111111111111101111111;
			22: value = 40'b1111111011111111111111111111111101111111;
			23: value = 40'b1111111011111111111111111111111101111111;
			24: value = 40'b1111111011111111111111111111111101111111;
			25: value = 40'b1111111011111111111111111111111101111111;
			26: value = 40'b1111111011111111111111111111111101111111;
			27: value = 40'b1111111011111111111111111111111101111111;
			28: value = 40'b1111111011111111111111111111111101111111;
			29: value = 40'b1111111011111111111111111111111101111111;
			30: value = 40'b1111111011111111111111111111111101111111;
			31: value = 40'b1111111011111111111111111111111101111111;
			32: value = 40'b1111100011111111111111111111111100011111;
			33: value = 40'b1111101111111111111111111111111111011111;
			34: value = 40'b1111101111111111111111111111111111011111;
			35: value = 40'b1111100000000000000000000000000000011111;
			36: value = 40'b1111111111111111111111111111111111111111;
			37: value = 40'b1111111111111111111111111111111111111111;
			38: value = 40'b1111111111111111111111111111111111111111;
			39: value = 40'b1111111111111111111111111111111111111111;
			default: value = 40'd0;
		endcase 

				
				end
				else begin
					case(row) //black square white rook
			0: value =  40'b0000000000000000000000000000000000000000;
			1: value =  40'b0000000000000000000000000000000000000000;
			2: value =  40'b0000000000000000000000000000000000000000;
			3: value =  40'b0000000000000000000000000000000000000000;
			4: value =  40'b0000000000000000000000000000000000000000;
			5: value =  40'b0000001111111000111111110001111111000000;
			6: value =  40'b0000001111111000111111110001111111000000;
			7: value =  40'b0000001111111000111111110001111111000000;
			8: value =  40'b0000001111111000111111110001111111000000;
			9: value=   40'b0000001111111111111111111111111111000000;
			10: value = 40'b0000001111111111111111111111111111000000;
			11: value = 40'b0000001111111111111111111111111111000000;
			12: value = 40'b0000001111111111111111111111111111000000;
			13: value = 40'b0000001111111111111111111111111111000000;
			14: value = 40'b0000001111111111111111111111111111000000;
			15: value = 40'b0000001111111111111111111111111111000000;
			16: value = 40'b0000000000001111111111111111000000000000;
			17: value = 40'b0000000000001111111111111111000000000000;
			18: value = 40'b0000000000001111111111111111000000000000;
			19: value = 40'b0000000000001111111111111111000000000000;
			20: value = 40'b0000000011111111111111111111111100000000;
			21: value = 40'b0000000011111111111111111111111100000000;
			22: value = 40'b0000000011111111111111111111111100000000;
			23: value = 40'b0000000011111111111111111111111100000000;
			24: value = 40'b0000000011111111111111111111111100000000;
			25: value = 40'b0000000011111111111111111111111100000000;
			26: value = 40'b0000000011111111111111111111111100000000;
			27: value = 40'b0000000011111111111111111111111100000000;
			28: value = 40'b0000000011111111111111111111111100000000;
			29: value = 40'b0000000011111111111111111111111100000000;
			30: value = 40'b0000000011111111111111111111111100000000;
			31: value = 40'b0000000011111111111111111111111100000000;
			32: value = 40'b0000000011111111111111111111111100000000;
			33: value = 40'b0000001111111111111111111111111111000000;
			34: value = 40'b0000001111111111111111111111111111000000;
			35: value = 40'b0000000000000000000000000000000000000000;
			36: value = 40'b0000000000000000000000000000000000000000;
			37: value = 40'b0000000000000000000000000000000000000000;
			38: value = 40'b0000000000000000000000000000000000000000;
			39: value = 40'b0000000000000000000000000000000000000000;
			default: value = 40'd0;
		endcase 
				end
			end
			else begin
				if(sqcolor)begin
						case(row)//white square black rook
			0: value =  40'b1111111111111111111111111111111111111111;
			1: value =  40'b1111111111111111111111111111111111111111;
			2: value =  40'b1111111111111111111111111111111111111111;
			3: value =  40'b1111111111111111111111111111111111111111;
			4: value =  40'b1111111111111111111111111111111111111111;
			5: value =  40'b1111110000000111000000001110000000111111;
			6: value =  40'b1111110000000111000000001110000000111111;
			7: value =  40'b1111110000000111000000001110000000111111;
			8: value =  40'b1111110000000111000000001110000000111111;
			9: value=   40'b1111110000000000000000000000000000111111;
			10: value = 40'b1111110000000000000000000000000000111111;
			11: value = 40'b1111110000000000000000000000000000111111;
			12: value = 40'b1111110000000000000000000000000000111111;
			13: value = 40'b1111110000000000000000000000000000111111;
			14: value = 40'b1111110000000000000000000000000000111111;
			15: value = 40'b1111110000000000000000000000000000111111;
			16: value = 40'b1111111111110000000000000000111111111111;
			17: value = 40'b1111111111110000000000000000111111111111;
			18: value = 40'b1111111111110000000000000000111111111111;
			19: value = 40'b1111111111110000000000000000111111111111;
			20: value = 40'b1111111100000000000000000000000011111111;
			21: value = 40'b1111111100000000000000000000000011111111;
			22: value = 40'b1111111100000000000000000000000011111111;
			23: value = 40'b1111111100000000000000000000000011111111;
			24: value = 40'b1111111100000000000000000000000011111111;
			25: value = 40'b1111111100000000000000000000000011111111;
			26: value = 40'b1111111100000000000000000000000011111111;
			27: value = 40'b1111111100000000000000000000000011111111;
			28: value = 40'b1111111100000000000000000000000011111111;
			29: value = 40'b1111111100000000000000000000000011111111;
			30: value = 40'b1111111100000000000000000000000011111111;
			31: value = 40'b1111111100000000000000000000000011111111;
			32: value = 40'b1111111100000000000000000000000011111111;
			33: value = 40'b1111110000000000000000000000000000111111;
			34: value = 40'b1111110000000000000000000000000000111111;
			35: value = 40'b1111111111111111111111111111111111111111;
			36: value = 40'b1111111111111111111111111111111111111111;
			37: value = 40'b1111111111111111111111111111111111111111;
			38: value = 40'b1111111111111111111111111111111111111111;
			39: value = 40'b1111111111111111111111111111111111111111;
			default: value = 40'd0;
		endcase 

				
				end
				else begin
						case(row) //black square black rook
			0: value =  40'b0000000000000000000000000000000000000000;
			1: value =  40'b0000000000000000000000000000000000000000;
			2: value =  40'b0000000000000000000000000000000000000000;
			3: value =  40'b0000000000000000000000000000000000000000;
			4: value =  40'b0000011111111101111111111011111111100000;
			5: value =  40'b0000010000000101000000001010000000100000;
			6: value =  40'b0000010000000101000000001010000000100000;
			7: value =  40'b0000010000000101000000001010000000100000;
			8: value =  40'b0000010000000111000000001110000000100000;
			9: value=   40'b0000010000000000000000000000000000100000;
			10: value = 40'b0000010000000000000000000000000000100000;
			11: value = 40'b0000010000000000000000000000000000100000;
			12: value = 40'b0000010000000000000000000000000000100000;
			13: value = 40'b0000010000000000000000000000000000100000;
			14: value = 40'b0000010000000000000000000000000000100000;
			15: value = 40'b0000010000000000000000000000000000100000;
			16: value = 40'b0000011111110000000000000000111111100000;
			17: value = 40'b0000000000010000000000000000100000000000;
			18: value = 40'b0000000000010000000000000000100000000000;
			19: value = 40'b0000000111110000000000000000111110000000;
			20: value = 40'b0000000100000000000000000000000010000000;
			21: value = 40'b0000000100000000000000000000000010000000;
			22: value = 40'b0000000100000000000000000000000010000000;
			23: value = 40'b0000000100000000000000000000000010000000;
			24: value = 40'b0000000100000000000000000000000010000000;
			25: value = 40'b0000000100000000000000000000000010000000;
			26: value = 40'b0000000100000000000000000000000010000000;
			27: value = 40'b0000000100000000000000000000000010000000;
			28: value = 40'b0000000100000000000000000000000010000000;
			29: value = 40'b0000000100000000000000000000000010000000;
			30: value = 40'b0000000100000000000000000000000010000000;
			31: value = 40'b0000000100000000000000000000000010000000;
			32: value = 40'b0000011100000000000000000000000011100000;
			33: value = 40'b0000010000000000000000000000000000100000;
			34: value = 40'b0000010000000000000000000000000000100000;
			35: value = 40'b0000011111111111111111111111111111100000;
			36: value = 40'b0000000000000000000000000000000000000000;
			37: value = 40'b0000000000000000000000000000000000000000;
			38: value = 40'b0000000000000000000000000000000000000000;
			39: value = 40'b0000000000000000000000000000000000000000;
			default: value = 40'd0;
		endcase 
				end
			end
		end
		
		
		horse:begin
			if(piece > 7)begin // if piece is white or black
				if(sqcolor)begin
						case(row)//white square white bishop
			0: value =  40'b1111111111111111111111111111111111111111;
			1: value =  40'b1111111111111111111111111111111111111111;
			2: value =  40'b1111111111111111111111111111111111111111;
			3: value =  40'b1111111111111111111111111111111111111111;
			4: value =  40'b1111111111111111100000000111111111111111;
			5: value =  40'b1111111111111111101111110111111111111111;
			6: value =  40'b1111111111111111011111111011111111111111;
			7: value =  40'b1111111111111110111111111101111111111111;
			8: value =  40'b1111111111111111011111111110111111111111;
			9: value =  40'b1111111111100000011111111110111111111111;
			10: value=  40'b1111111111101111111111111111011111111111;
			11: value = 40'b1111111111011111111111111111011111111111;
			12: value = 40'b1111111110111111111111111110111111111111;
			13: value = 40'b1111111101111111111111111101111111111111;
			14: value = 40'b1111111101111111111111111101111111111111;
			15: value = 40'b1111111101111111111111111101111111111111;
			16: value = 40'b1111111101111110011111111101111111111111;
			17: value = 40'b1111111101111101011111111101111111111111;
			18: value = 40'b1111111101111011011111111101111111111111;
			19: value = 40'b1111111100000001111111111101111111111111;
			20: value = 40'b1111111111111101111111111101111111111111;
			21: value = 40'b1111111111110001111111111101111111111111;
			22: value = 40'b1111111111110111111111111101111111111111;
			23: value = 40'b1111111111110111111111111101111111111111;
			24: value = 40'b1111111111110111111111111101111111111111;
			25: value = 40'b1111111111101111111111111101111111111111;
			26: value = 40'b1111111111101111111111111101111111111111;
			27: value = 40'b1111111111101111111111111101111111111111;
			28: value = 40'b1111111111011111111111111110111111111111;
			29: value = 40'b1111111111011111111111111110111111111111;
			30: value = 40'b1111111100011111111111111110001111111111;
			31: value = 40'b1111000001111111111111111111100000111111;
			32: value = 40'b1111011111111111111111111111111110111111;
			33: value = 40'b1111011111111111111111111111111110111111;
			34: value = 40'b1111011111111111111111111111111110111111;
			35: value = 40'b1111000000000000000000000000000000111111;
			36: value = 40'b1111111111111111111111111111111111111111;
			37: value = 40'b1111111111111111111111111111111111111111;
			38: value = 40'b1111111111111111111111111111111111111111;
			39: value = 40'b1111111111111111111111111111111111111111;
			default: value = 40'd0;
		endcase 
				
				end
				else begin
					case(row) //black square white bishop
			0: value =  40'b0000000000000000000000000000000000000000;
			1: value =  40'b0000000000000000000000000000000000000000;
			2: value =  40'b0000000000000000000000000000000000000000;
			3: value =  40'b0000000000000000000000000000000000000000;
			4: value =  40'b0000000000000000000000000000000000000000;
			5: value =  40'b0000000000000000001111110000000000000000;
			6: value =  40'b0000000000000000011111111000000000000000;
			7: value =  40'b0000000000000000111111111100000000000000;
			8: value =  40'b0000000000000000011111111110000000000000;
			9: value =  40'b0000000000000100011111111110000000000000;
			10: value=  40'b0000000000001111111111111111000000000000;
			11: value = 40'b0000000000011111111111111111000000000000;
			12: value = 40'b0000000000111111111111111110000000000000;
			13: value = 40'b0000000001111111111111111100000000000000;
			14: value = 40'b0000000001111111111111111100000000000000;
			15: value = 40'b0000000001111111111111111100000000000000;
			16: value = 40'b0000000001111110011111111100000000000000;
			17: value = 40'b0000000001111100011111111100000000000000;
			18: value = 40'b0000000001111000011111111100000000000000;
			19: value = 40'b0000000000000001111111111100000000000000;
			20: value = 40'b0000000000000001111111111100000000000000;
			21: value = 40'b0000000000000001111111111100000000000000;
			22: value = 40'b0000000000000111111111111100000000000000;
			23: value = 40'b0000000000000111111111111100000000000000;
			24: value = 40'b0000000000000111111111111100000000000000;
			25: value = 40'b0000000000001111111111111100000000000000;
			26: value = 40'b0000000000001111111111111100000000000000;
			27: value = 40'b0000000000001111111111111100000000000000;
			28: value = 40'b0000000000011111111111111110000000000000;
			29: value = 40'b0000000000011111111111111110000000000000;
			30: value = 40'b0000000000011111111111111110000000000000;
			31: value = 40'b0000000001111111111111111111100000000000;
			32: value = 40'b0000011111111111111111111111111110000000;
			33: value = 40'b0000011111111111111111111111111110000000;
			34: value = 40'b0000011111111111111111111111111110000000;
			35: value = 40'b0000000000000000000000000000000000000000;
			36: value = 40'b0000000000000000000000000000000000000000;
			37: value = 40'b0000000000000000000000000000000000000000;
			38: value = 40'b0000000000000000000000000000000000000000;
			39: value = 40'b0000000000000000000000000000000000000000;
			default: value = 40'd0;
		endcase 

				end
			end
			else begin
				if(sqcolor)begin
				case(row)//white square black bishop
			0: value =  40'b1111111111111111111111111111111111111111;
			1: value =  40'b1111111111111111111111111111111111111111;
			2: value =  40'b1111111111111111111111111111111111111111;
			3: value =  40'b1111111111111111111111111111111111111111;
			4: value =  40'b1111111111111111111111111111111111111111;
			5: value =  40'b1111111111111111110000001111111111111111;
			6: value =  40'b1111111111111111100000000111111111111111;
			7: value =  40'b1111111111111111000000000011111111111111;
			8: value =  40'b1111111111111111100000000001111111111111;
			9: value =  40'b1111111111111011100000000001111111111111;
			10: value=  40'b1111111111110000000000000000111111111111;
			11: value = 40'b1111111111100000000000000000111111111111;
			12: value = 40'b1111111111000000000000000001111111111111;
			13: value = 40'b1111111110000000000000000011111111111111;
			14: value = 40'b1111111110000000000000000011111111111111;
			15: value = 40'b1111111110000000000000000011111111111111;
			16: value = 40'b1111111110000001100000000011111111111111;
			17: value = 40'b1111111110000011100000000011111111111111;
			18: value = 40'b1111111110000111100000000011111111111111;
			19: value = 40'b1111111111111110000000000011111111111111;
			20: value = 40'b1111111111111110000000000011111111111111;
			21: value = 40'b1111111111111110000000000011111111111111;
			22: value = 40'b1111111111111000000000000011111111111111;
			23: value = 40'b1111111111111000000000000011111111111111;
			24: value = 40'b1111111111111000000000000011111111111111;
			25: value = 40'b1111111111110000000000000011111111111111;
			26: value = 40'b1111111111110000000000000011111111111111;
			27: value = 40'b1111111111110000000000000011111111111111;
			28: value = 40'b1111111111100000000000000001111111111111;
			29: value = 40'b1111111111100000000000000001111111111111;
			30: value = 40'b1111111111100000000000000001111111111111;
			31: value = 40'b1111111110000000000000000000011111111111;
			32: value = 40'b1111100000000000000000000000000001111111;
			33: value = 40'b1111100000000000000000000000000001111111;
			34: value = 40'b1111100000000000000000000000000001111111;
			35: value = 40'b1111111111111111111111111111111111111111;
			36: value = 40'b1111111111111111111111111111111111111111;
			37: value = 40'b1111111111111111111111111111111111111111;
			38: value = 40'b1111111111111111111111111111111111111111;
			39: value = 40'b1111111111111111111111111111111111111111;
			default: value = 40'd0;
		endcase 	
				
				end
				else begin
						case(row) //black square black bishop
			0: value =  40'b0000000000000000000000000000000000000000;
			1: value =  40'b0000000000000000000000000000000000000000;
			2: value =  40'b0000000000000000000000000000000000000000;
			3: value =  40'b0000000000000000000000000000000000000000;
			4: value =  40'b0000000000000000011111111000000000000000;
			5: value =  40'b0000000000000000010000001000000000000000;
			6: value =  40'b0000000000000000100000000100000000000000;
			7: value =  40'b0000000000000001000000000010000000000000;
			8: value =  40'b0000000000000000100000000001000000000000;
			9: value =  40'b0000000000011111100000000001000000000000;
			10: value=  40'b0000000000010000000000000000100000000000;
			11: value = 40'b0000000000100000000000000000100000000000;
			12: value = 40'b0000000001000000000000000001000000000000;
			13: value = 40'b0000000010000000000000000010000000000000;
			14: value = 40'b0000000010000000000000000010000000000000;
			15: value = 40'b0000000010000000000000000010000000000000;
			16: value = 40'b0000000010000001100000000010000000000000;
			17: value = 40'b0000000010000010100000000010000000000000;
			18: value = 40'b0000000010000100100000000010000000000000;
			19: value = 40'b0000000011111110000000000010000000000000;
			20: value = 40'b0000000000000010000000000010000000000000;
			21: value = 40'b0000000000001110000000000010000000000000;
			22: value = 40'b0000000000001000000000000010000000000000;
			23: value = 40'b0000000000001000000000000010000000000000;
			24: value = 40'b0000000000001000000000000010000000000000;
			25: value = 40'b0000000000010000000000000010000000000000;
			26: value = 40'b0000000000010000000000000010000000000000;
			27: value = 40'b0000000000010000000000000010000000000000;
			28: value = 40'b0000000000100000000000000001000000000000;
			29: value = 40'b0000000000100000000000000001000000000000;
			30: value = 40'b0000000011100000000000000001110000000000;
			31: value = 40'b0000111110000000000000000000011111000000;
			32: value = 40'b0000100000000000000000000000000001000000;
			33: value = 40'b0000100000000000000000000000000001000000;
			34: value = 40'b0000100000000000000000000000000001000000;
			35: value = 40'b0000111111111111111111111111111111000000;
			36: value = 40'b0000000000000000000000000000000000000000;
			37: value = 40'b0000000000000000000000000000000000000000;
			38: value = 40'b0000000000000000000000000000000000000000;
			39: value = 40'b0000000000000000000000000000000000000000;
			default: value = 40'd0;
		endcase

				end
			end
		end
		
		bishop:begin
			if(piece > 7)begin // if piece is white or black
				if(sqcolor)begin
					case(row)//white square white bishop
			0: value =  40'b1111111111111111111111111111111111111111;
			1: value =  40'b1111111111111111111111111111111111111111;
			2: value =  40'b1111111111111111111111111111111111111111;
			3: value =  40'b1111111111111111111111111111111111111111;
			4: value =  40'b1111111111111111100000011111111111111111;
			5: value =  40'b1111111111111111101111011111111111111111;
			6: value =  40'b1111111111111111101111011111111111111111;
			7: value =  40'b1111111111111111101111011111111111111111;
			8: value =  40'b1111111111111111100110011111111111111111;
			9: value =  40'b1111111111111111101111011111111111111111;
			10: value=  40'b1111111111111111110111101111111111111111;
			11: value = 40'b1111111111111111001011110111111111111111;
			12: value = 40'b1111111111111110110101111011111111111111;
			13: value = 40'b1111111111111101111010111101111111111111;
			14: value = 40'b1111111111111011111100111110111111111111;
			15: value = 40'b1111111111110111111111111111011111111111;
			16: value = 40'b1111111111101111111111111111101111111111;
			17: value = 40'b1111111111011111111111111111110111111111;
			18: value = 40'b1111111110111111111111111111111011111111;
			19: value = 40'b1111111101111111111111111111111101111111;
			20: value = 40'b1111111011111111111111111111111110111111;
			21: value = 40'b1111110111111111111111111111111111011111;
			22: value = 40'b1111110111111111111111111111111111011111;
			23: value = 40'b1111110111111111111111111111111111011111;
			24: value = 40'b1111110111111111111111111111111111011111;
			25: value = 40'b1111110111111111111111111111111111011111;
			26: value = 40'b1111110111111111111111111111111111011111;
			27: value = 40'b1111110111111111111111111111111111011111;
			28: value = 40'b1111111011111111111111111111111110111111;
			29: value = 40'b1111111101111111111111111111111101111111;
			30: value = 40'b1111111110111111111111111111111011111111;
			31: value = 40'b1111111000001111111111111111110000011111;
			32: value = 40'b1111111011111111111111111111111111011111;
			33: value = 40'b1111111011111111111111111111111111011111;
			34: value = 40'b1111111011111111111111111111111111011111;
			35: value = 40'b1111111000000000000000000000000000011111;
			36: value = 40'b1111111111111111111111111111111111111111;
			37: value = 40'b1111111111111111111111111111111111111111;
			38: value = 40'b1111111111111111111111111111111111111111;
			39: value = 40'b1111111111111111111111111111111111111111;
			default: value = 40'd0;
		endcase 
				
				end
				else begin
					case(row) //black square white bishop
			0: value =  40'b0000000000000000000000000000000000000000;
			1: value =  40'b0000000000000000000000000000000000000000;
			2: value =  40'b0000000000000000000000000000000000000000;
			3: value =  40'b0000000000000000000000000000000000000000;
			4: value =  40'b0000000000000000000000000000000000000000;
			5: value =  40'b0000000000000000001111000000000000000000;
			6: value =  40'b0000000000000000001111000000000000000000;
			7: value =  40'b0000000000000000001111000000000000000000;
			8: value =  40'b0000000000000000000110000000000000000000;
			9: value =  40'b0000000000000000001111000000000000000000;
			10: value=  40'b0000000000000000000111100000000000000000;
			11: value = 40'b0000000000000000000011110000000000000000;
			12: value = 40'b0000000000000000110001111000000000000000;
			13: value = 40'b0000000000000001111000111100000000000000;
			14: value = 40'b0000000000000011111100111110000000000000;
			15: value = 40'b0000000000000111111111111111000000000000;
			16: value = 40'b0000000000001111111111111111100000000000;
			17: value = 40'b0000000000011111111111111111110000000000;
			18: value = 40'b0000000000111111111111111111111000000000;
			19: value = 40'b0000000001111111111111111111111100000000;
			20: value = 40'b0000000011111111111111111111111110000000;
			21: value = 40'b0000000111111111111111111111111111000000;
			22: value = 40'b0000000111111111111111111111111111000000;
			23: value = 40'b0000000111111111111111111111111111000000;
			24: value = 40'b0000000111111111111111111111111111000000;
			25: value = 40'b0000000111111111111111111111111111000000;
			26: value = 40'b0000000111111111111111111111111111000000;
			27: value = 40'b0000000111111111111111111111111111000000;
			28: value = 40'b0000000011111111111111111111111110000000;
			29: value = 40'b0000000001111111111111111111111100000000;
			30: value = 40'b0000000000111111111111111111111000000000;
			31: value = 40'b0000000000001111111111111111110000000000;
			32: value = 40'b0000000011111111111111111111111111000000;
			33: value = 40'b0000000011111111111111111111111111000000;
			34: value = 40'b0000000011111111111111111111111111000000;
			35: value = 40'b0000000000000000000000000000000000000000;
			36: value = 40'b0000000000000000000000000000000000000000;
			37: value = 40'b0000000000000000000000000000000000000000;
			38: value = 40'b0000000000000000000000000000000000000000;
			39: value = 40'b0000000000000000000000000000000000000000;
			default: value = 40'd0;
		endcase 
				end
			end
			else begin
				if(sqcolor)begin
						case(row)//white square black bishop
			0: value =  40'b1111111111111111111111111111111111111111;
			1: value =  40'b1111111111111111111111111111111111111111;
			2: value =  40'b1111111111111111111111111111111111111111;
			3: value =  40'b1111111111111111111111111111111111111111;
			4: value =  40'b1111111111111111111111111111111111111111;
			5: value =  40'b1111111111111111110000111111111111111111;
			6: value =  40'b1111111111111111110000111111111111111111;
			7: value =  40'b1111111111111111110000111111111111111111;
			8: value =  40'b1111111111111111111001111111111111111111;
			9: value =  40'b1111111111111111110000111111111111111111;
			10: value=  40'b1111111111111111111000011111111111111111;
			11: value = 40'b1111111111111111111100001111111111111111;
			12: value = 40'b1111111111111111001110000111111111111111;
			13: value = 40'b1111111111111110000111000011111111111111;
			14: value = 40'b1111111111111100000011000001111111111111;
			15: value = 40'b1111111111111000000000000000111111111111;
			16: value = 40'b1111111111110000000000000000011111111111;
			17: value = 40'b1111111111100000000000000000001111111111;
			18: value = 40'b1111111111000000000000000000000111111111;
			19: value = 40'b1111111110000000000000000000000011111111;
			20: value = 40'b1111111100000000000000000000000001111111;
			21: value = 40'b1111111000000000000000000000000000111111;
			22: value = 40'b1111111000000000000000000000000000111111;
			23: value = 40'b1111111000000000000000000000000000111111;
			24: value = 40'b1111111000000000000000000000000000111111;
			25: value = 40'b1111111000000000000000000000000000111111;
			26: value = 40'b1111111000000000000000000000000000111111;
			27: value = 40'b1111111000000000000000000000000000111111;
			28: value = 40'b1111111100000000000000000000000001111111;
			29: value = 40'b1111111110000000000000000000000011111111;
			30: value = 40'b1111111111000000000000000000000111111111;
			31: value = 40'b1111111111110000000000000000001111111111;
			32: value = 40'b1111111100000000000000000000000000111111;
			33: value = 40'b1111111100000000000000000000000000111111;
			34: value = 40'b1111111100000000000000000000000000111111;
			35: value = 40'b1111111111111111111111111111111111111111;
			36: value = 40'b1111111111111111111111111111111111111111;
			37: value = 40'b1111111111111111111111111111111111111111;
			38: value = 40'b1111111111111111111111111111111111111111;
			39: value = 40'b1111111111111111111111111111111111111111;
			default: value = 40'd0;
		endcase 
				
				end
				else begin
					case(row) //black square black bishop
			0: value =  40'b0000000000000000000000000000000000000000;
			1: value =  40'b0000000000000000000000000000000000000000;
			2: value =  40'b0000000000000000000000000000000000000000;
			3: value =  40'b0000000000000000000000000000000000000000;
			4: value =  40'b0000000000000000011111100000000000000000;
			5: value =  40'b0000000000000000010000100000000000000000;
			6: value =  40'b0000000000000000010000100000000000000000;
			7: value =  40'b0000000000000000010000100000000000000000;
			8: value =  40'b0000000000000000011001100000000000000000;
			9: value =  40'b0000000000000000010000100000000000000000;
			10: value=  40'b0000000000000000001000010000000000000000;
			11: value = 40'b0000000000000000110100001000000000000000;
			12: value = 40'b0000000000000001001010000100000000000000;
			13: value = 40'b0000000000000010000101000010000000000000;
			14: value = 40'b0000000000000100000011000001000000000000;
			15: value = 40'b0000000000001000000000000000100000000000;
			16: value = 40'b0000000000010000000000000000010000000000;
			17: value = 40'b0000000000100000000000000000001000000000;
			18: value = 40'b0000000001000000000000000000000100000000;
			19: value = 40'b0000000010000000000000000000000010000000;
			20: value = 40'b0000000100000000000000000000000001000000;
			21: value = 40'b0000001000000000000000000000000000100000;
			22: value = 40'b0000001000000000000000000000000000100000;
			23: value = 40'b0000001000000000000000000000000000100000;
			24: value = 40'b0000001000000000000000000000000000100000;
			25: value = 40'b0000001000000000000000000000000000100000;
			26: value = 40'b0000001000000000000000000000000000100000;
			27: value = 40'b0000001000000000000000000000000000100000;
			28: value = 40'b0000000100000000000000000000000001000000;
			29: value = 40'b0000000010000000000000000000000010000000;
			30: value = 40'b0000000001000000000000000000000100000000;
			31: value = 40'b0000000111110000000000000000001111100000;
			32: value = 40'b0000000100000000000000000000000000100000;
			33: value = 40'b0000000100000000000000000000000000100000;
			34: value = 40'b0000000100000000000000000000000000100000;
			35: value = 40'b0000000111111111111111111111111111100000;
			36: value = 40'b0000000000000000000000000000000000000000;
			37: value = 40'b0000000000000000000000000000000000000000;
			38: value = 40'b0000000000000000000000000000000000000000;
			39: value = 40'b0000000000000000000000000000000000000000;
			default: value = 40'd0;
		endcase 
				end
			end
		end
		
		queen:begin
			if(piece > 7)begin // if piece is white or black
				if(sqcolor)begin
					case(row)//white square white queen
			0: value =  40'b1111111111111111111111111111111111111111;
			1: value =  40'b1111111111111111111111111111111111111111;
			2: value =  40'b1111111111111111111111111111111111111111;
			3: value =  40'b1111111111111111111111111111111111111111;
			4: value =  40'b1111111111111111111001111111111111111111;
			5: value =  40'b1111111111111111110110111111111111111111;
			6: value =  40'b1111111111111111101111011111111111111111;
			7: value =  40'b1111111111111111011111101111111111111111;
			8: value =  40'b1111111111111110111111110111111111111111;
			9: value =  40'b1111111111111110111111110111111111111111;
			10: value=  40'b1111111111111111011111101111111111111111;
			11: value = 40'b1111111111111111101111011111111111111111;
			12: value = 40'b1111111111111111000110001111111111111111;
			13: value = 40'b1111111111111100011111100011111111111111;
			14: value = 40'b1111111100000001111111111000000011111111;
			15: value = 40'b1111111101100111111111111110011011111111;
			16: value = 40'b1111111101111111111111111111111011111111;
			17: value = 40'b1111111101111111111111111111111011111111;
			18: value = 40'b1111111101111111111111111111111011111111;
			19: value = 40'b1111111101111111111111111111111011111111;
			20: value = 40'b1111111101111111111111111111111011111111;
			21: value = 40'b1111111100011111111111111111100011111111;
			22: value = 40'b1111111111100000111111110000011111111111;
			23: value = 40'b1111111111111110111111110111111111111111;
			24: value = 40'b1111111111111110111111110111111111111111;
			25: value = 40'b1111111111111110111111110111111111111111;
			26: value = 40'b1111111111111110111111110111111111111111;
			27: value = 40'b1111111111111110111111110111111111111111;
			28: value = 40'b1111111111111000111111110001111111111111;
			29: value = 40'b1111111111111011111111111101111111111111;
			30: value = 40'b1111111110000011111111111100000111111111;
			31: value = 40'b1111111110111111111111111111110111111111;
			32: value = 40'b1111111110111111111111111111110111111111;
			33: value = 40'b1111111110111111111111111111110111111111;
			34: value = 40'b1111111110111111111111111111110111111111;
			35: value = 40'b1111111110000000000000000000000111111111;
			36: value = 40'b1111111111111111111111111111111111111111;
			37: value = 40'b1111111111111111111111111111111111111111;
			38: value = 40'b1111111111111111111111111111111111111111;
			39: value = 40'b1111111111111111111111111111111111111111;
			default: value = 40'd0;
		endcase
				
				end
				else begin
					case(row) //black square white queen
			0: value =  40'b0000000000000000000000000000000000000000;
			1: value =  40'b0000000000000000000000000000000000000000;
			2: value =  40'b0000000000000000000000000000000000000000;
			3: value =  40'b0000000000000000000000000000000000000000;
			4: value =  40'b0000000000000000000000000000000000000000;
			5: value =  40'b0000000000000000000110000000000000000000;
			6: value =  40'b0000000000000000001111000000000000000000;
			7: value =  40'b0000000000000000011111100000000000000000;
			8: value =  40'b0000000000000000111111110000000000000000;
			9: value =  40'b0000000000000000111111110000000000000000;
			10: value=  40'b0000000000000000011111100000000000000000;
			11: value = 40'b0000000000000000001111000000000000000000;
			12: value = 40'b0000000000000000000110000000000000000000;
			13: value = 40'b0000000000000000011111100000000000000000;
			14: value = 40'b0000000000000001111111111000000000000000;
			15: value = 40'b0000000001100111111111111110011000000000;
			16: value = 40'b0000000001111111111111111111111000000000;
			17: value = 40'b0000000001111111111111111111111000000000;
			18: value = 40'b0000000001111111111111111111111000000000;
			19: value = 40'b0000000001111111111111111111111000000000;
			20: value = 40'b0000000000111111111111111111110000000000;
			21: value = 40'b0000000000011111111111111111100000000000;
			22: value = 40'b0000000000000000111111110000000000000000;
			23: value = 40'b0000000000000000111111110000000000000000;
			24: value = 40'b0000000000000000111111110000000000000000;
			25: value = 40'b0000000000000000111111110000000000000000;
			26: value = 40'b0000000000000000111111110000000000000000;
			27: value = 40'b0000000000000000111111110000000000000000;
			28: value = 40'b0000000000000000111111110000000000000000;
			29: value = 40'b0000000000000011111111111100000000000000;
			30: value = 40'b0000000000000011111111111100000000000000;
			31: value = 40'b0000000000111111111111111111110000000000;
			32: value = 40'b0000000000111111111111111111110000000000;
			33: value = 40'b0000000000111111111111111111110000000000;
			34: value = 40'b0000000000111111111111111111110000000000;
			35: value = 40'b0000000000000000000000000000000000000000;
			36: value = 40'b0000000000000000000000000000000000000000;
			37: value = 40'b0000000000000000000000000000000000000000;
			38: value = 40'b0000000000000000000000000000000000000000;
			39: value = 40'b0000000000000000000000000000000000000000;
			default: value = 40'd0;
		endcase 
				end
			end
			else begin
				if(sqcolor)begin
				case(row)//white square black queen
			0: value =  40'b1111111111111111111111111111111111111111;
			1: value =  40'b1111111111111111111111111111111111111111;
			2: value =  40'b1111111111111111111111111111111111111111;
			3: value =  40'b1111111111111111111111111111111111111111;
			4: value =  40'b1111111111111111111111111111111111111111;
			5: value =  40'b1111111111111111111001111111111111111111;
			6: value =  40'b1111111111111111110000111111111111111111;
			7: value =  40'b1111111111111111100000011111111111111111;
			8: value =  40'b1111111111111111000000001111111111111111;
			9: value =  40'b1111111111111111000000001111111111111111;
			10: value=  40'b1111111111111111100000011111111111111111;
			11: value = 40'b1111111111111111110000111111111111111111;
			12: value = 40'b1111111111111111111001111111111111111111;
			13: value = 40'b1111111111111111100000011111111111111111;
			14: value = 40'b1111111111111110000000000111111111111111;
			15: value = 40'b1111111110011000000000000001100111111111;
			16: value = 40'b1111111110000000000000000000000111111111;
			17: value = 40'b1111111110000000000000000000000111111111;
			18: value = 40'b1111111110000000000000000000000111111111;
			19: value = 40'b1111111110000000000000000000000111111111;
			20: value = 40'b1111111111000000000000000000001111111111;
			21: value = 40'b1111111111100000000000000000011111111111;
			22: value = 40'b1111111111110000000000000000111111111111;
			23: value = 40'b1111111111111111000000001111111111111111;
			24: value = 40'b1111111111111111000000001111111111111111;
			25: value = 40'b1111111111111111000000001111111111111111;
			26: value = 40'b1111111111111111000000001111111111111111;
			27: value = 40'b1111111111111111000000001111111111111111;
			28: value = 40'b1111111111111111000000001111111111111111;
			29: value = 40'b1111111111111100000000000011111111111111;
			30: value = 40'b1111111111111100000000000011111111111111;
			31: value = 40'b1111111111000000000000000000001111111111;
			32: value = 40'b1111111111000000000000000000001111111111;
			33: value = 40'b1111111111000000000000000000001111111111;
			34: value = 40'b1111111111000000000000000000001111111111;
			35: value = 40'b1111111111111111111111111111111111111111;
			36: value = 40'b1111111111111111111111111111111111111111;
			37: value = 40'b1111111111111111111111111111111111111111;
			38: value = 40'b1111111111111111111111111111111111111111;
			39: value = 40'b1111111111111111111111111111111111111111;
			default: value = 40'd0;
		endcase
				
				end
				else begin
						case(row) //black square black queen
			0: value =  40'b0000000000000000000000000000000000000000;
			1: value =  40'b0000000000000000000000000000000000000000;
			2: value =  40'b0000000000000000000000000000000000000000;
			3: value =  40'b0000000000000000000000000000000000000000;
			4: value =  40'b0000000000000000000110000000000000000000;
			5: value =  40'b0000000000000000001001000000000000000000;
			6: value =  40'b0000000000000000010000100000000000000000;
			7: value =  40'b0000000000000000100000010000000000000000;
			8: value =  40'b0000000000000001000000001000000000000000;
			9: value =  40'b0000000000000001000000001000000000000000;
			10: value=  40'b0000000000000000100000010000000000000000;
			11: value = 40'b0000000000000000010000100000000000000000;
			12: value = 40'b0000000000000000111001110000000000000000;
			13: value = 40'b0000000000000011100000011100000000000000;
			14: value = 40'b0000000011111110000000000111111100000000;
			15: value = 40'b0000000010011000000000000001100100000000;
			16: value = 40'b0000000010000000000000000000000100000000;
			17: value = 40'b0000000010000000000000000000000100000000;
			18: value = 40'b0000000010000000000000000000000100000000;
			19: value = 40'b0000000010000000000000000000000100000000;
			20: value = 40'b0000000010000000000000000000000100000000;
			21: value = 40'b0000000011100000000000000000011100000000;
			22: value = 40'b0000000000011111000000001111100000000000;
			23: value = 40'b0000000000000001000000001000000000000000;
			24: value = 40'b0000000000000001000000001000000000000000;
			25: value = 40'b0000000000000001000000001000000000000000;
			26: value = 40'b0000000000000001000000001000000000000000;
			27: value = 40'b0000000000000001000000001000000000000000;
			28: value = 40'b0000000000000111000000001110000000000000;
			29: value = 40'b0000000000000100000000000010000000000000;
			30: value = 40'b0000000001111100000000000011111000000000;
			31: value = 40'b0000000001000000000000000000001000000000;
			32: value = 40'b0000000001000000000000000000001000000000;
			33: value = 40'b0000000001000000000000000000001000000000;
			34: value = 40'b0000000001000000000000000000001000000000;
			35: value = 40'b0000000001111111111111111111111000000000;
			36: value = 40'b0000000000000000000000000000000000000000;
			37: value = 40'b0000000000000000000000000000000000000000;
			38: value = 40'b0000000000000000000000000000000000000000;
			39: value = 40'b0000000000000000000000000000000000000000;
			default: value = 40'd0;
		endcase 
				end
			end
		end
		
		king:begin
			if(piece > 7)begin // if piece is white or black
				if(sqcolor)begin
				 case(row)//white square white king
					0: value =  40'b1111111111111111111111111111111111111111;
					1: value =  40'b1111111111111111111111111111111111111111;
					2: value =  40'b1111111111111111111111111111111111111111;
					3: value =  40'b1111111111111111111111111111111111111111;
					4: value =  40'b1111111111111111111001111111111111111111;
					5: value =  40'b1111111111111111110110111111111111111111;
					6: value =  40'b1111111111111111000110001111111111111111;
					7: value =  40'b1111111111111111011111101111111111111111;
					8: value =  40'b1111111111111111000110001111111111111111;
					9: value=   40'b1111111111111111110110111111111111111111;
					10: value = 40'b1111111111111111110110111111111111111111;
					11: value = 40'b1111111111111111101111011111111111111111;
					12: value = 40'b1111111111111111011111101111111111111111;
					13: value = 40'b1111111111111110111111110111111111111111;
					14: value = 40'b1111111111111101111111111011111111111111;
					15: value = 40'b1111111111111011111111111101111111111111;
					16: value = 40'b1111111111111011111111111101111111111111;
					17: value = 40'b1111111111111101111111111011111111111111;
					18: value = 40'b1111111111111110111111110111111111111111;
					19: value = 40'b1111111111111111011111101111111111111111;
					20: value = 40'b1111111111111000001111000001111111111111;
					21: value = 40'b1111111111111011111111111101111111111111;
					22: value = 40'b1111111111111011111111111101111111111111;
					23: value = 40'b1111111111111000001111000001111111111111;
					24: value = 40'b1111111111111111101111011111111111111111;
					25: value = 40'b1111111111111111011111101111111111111111;
					26: value = 40'b1111111111111111011111101111111111111111;
					27: value = 40'b1111111111111110111111110111111111111111;
					28: value = 40'b1111111111111110111111110111111111111111;
					29: value = 40'b1111111111111101111111111011111111111111;
					30: value = 40'b1111111111111101111111111011111111111111;
					31: value = 40'b1111111111111011111111111101111111111111;
					32: value = 40'b1111111111000011111111111100001111111111;
					33: value = 40'b1111111111011111111111111111101111111111;
					34: value = 40'b1111111111011111111111111111101111111111;
					35: value = 40'b1111111111000000000000000000001111111111;
					36: value = 40'b1111111111111111111111111111111111111111;
					37: value = 40'b1111111111111111111111111111111111111111;
					38: value = 40'b1111111111111111111111111111111111111111;
					39: value = 40'b1111111111111111111111111111111111111111;
					default: value = 40'd0;
			  endcase
				
				end
				else begin
					case(row)//black square white king
						0: value =  40'b0000000000000000000000000000000000000000;
						1: value =  40'b0000000000000000000000000000000000000000;
						2: value =  40'b0000000000000000000000000000000000000000;
						3: value =  40'b0000000000000000000000000000000000000000;
						4: value =  40'b0000000000000000000000000000000000000000;
						5: value =  40'b0000000000000000000110000000000000000000;
						6: value =  40'b0000000000000000000110000000000000000000;
						7: value =  40'b0000000000000000011111100000000000000000;
						8: value =  40'b0000000000000000000110000000000000000000;
						9: value=   40'b0000000000000000000110000000000000000000;
						10: value = 40'b0000000000000000000110000000000000000000;
						11: value = 40'b0000000000000000001111000000000000000000;
						12: value = 40'b0000000000000000011111100000000000000000;
						13: value = 40'b0000000000000000111111110000000000000000;
						14: value = 40'b0000000000000001111111111000000000000000;
						15: value = 40'b0000000000000011111111111100000000000000;
						16: value = 40'b0000000000000011111111111100000000000000;
						17: value = 40'b0000000000000001111111111000000000000000;
						18: value = 40'b0000000000000000111111110000000000000000;
						19: value = 40'b0000000000000000011111100000000000000000;
						20: value = 40'b0000000000000000001111000000000000000000;
						21: value = 40'b0000000000000011111111111100000000000000;
						22: value = 40'b0000000000000011111111111100000000000000;
						23: value = 40'b0000000000000000001111000000000000000000;
						24: value = 40'b0000000000000000001111000000000000000000;
						25: value = 40'b0000000000000000011111100000000000000000;
						26: value = 40'b0000000000000000011111100000000000000000;
						27: value = 40'b0000000000000000111111110000000000000000;
						28: value = 40'b0000000000000000111111110000000000000000;
						29: value = 40'b0000000000000001111111111000000000000000;
						30: value = 40'b0000000000000001111111111000000000000000;
						31: value = 40'b0000000000000011111111111100000000000000;
						32: value = 40'b0000000000000011111111111100000000000000;
						33: value = 40'b0000000000011111111111111111100000000000;
						34: value = 40'b0000000000011111111111111111100000000000;
						35: value = 40'b0000000000000000000000000000000000000000;
						36: value = 40'b0000000000000000000000000000000000000000;
						37: value = 40'b0000000000000000000000000000000000000000;
						38: value = 40'b0000000000000000000000000000000000000000;
						39: value = 40'b0000000000000000000000000000000000000000;
						default: value = 40'd0;
				  endcase
							end
			end
			else begin
				if(sqcolor)begin
					case(row)//white square black king
						0: value =  40'b1111111111111111111111111111111111111111;
						1: value =  40'b1111111111111111111111111111111111111111;
						2: value =  40'b1111111111111111111111111111111111111111;
						3: value =  40'b1111111111111111111111111111111111111111;
						4: value =  40'b1111111111111111111111111111111111111111;
						5: value =  40'b1111111111111111111001111111111111111111;
						6: value =  40'b1111111111111111111001111111111111111111;
						7: value =  40'b1111111111111111100000011111111111111111;
						8: value =  40'b1111111111111111111001111111111111111111;
						9: value=   40'b1111111111111111111001111111111111111111;
						10: value = 40'b1111111111111111111001111111111111111111;
						11: value = 40'b1111111111111111110000111111111111111111;
						12: value = 40'b1111111111111111100000011111111111111111;
						13: value = 40'b1111111111111111000000001111111111111111;
						14: value = 40'b1111111111111110000000000111111111111111;
						15: value = 40'b1111111111111100000000000011111111111111;
						16: value = 40'b1111111111111100000000000011111111111111;
						17: value = 40'b1111111111111110000000000111111111111111;
						18: value = 40'b1111111111111111000000001111111111111111;
						19: value = 40'b1111111111111111100000011111111111111111;
						20: value = 40'b1111111111111111110000111111111111111111;
						21: value = 40'b1111111111111100000000000011111111111111;
						22: value = 40'b1111111111111100000000000011111111111111;
						23: value = 40'b1111111111111111110000111111111111111111;
						24: value = 40'b1111111111111111110000111111111111111111;
						25: value = 40'b1111111111111111100000011111111111111111;
						26: value = 40'b1111111111111111100000011111111111111111;
						27: value = 40'b1111111111111111000000001111111111111111;
						28: value = 40'b1111111111111111000000001111111111111111;
						29: value = 40'b1111111111111110000000000111111111111111;
						30: value = 40'b1111111111111110000000000111111111111111;
						31: value = 40'b1111111111111100000000000011111111111111;
						32: value = 40'b1111111111111100000000000011111111111111;
						33: value = 40'b1111111111100000000000000000011111111111;
						34: value = 40'b1111111111100000000000000000011111111111;
						35: value = 40'b1111111111111111111111111111111111111111;
						36: value = 40'b1111111111111111111111111111111111111111;
						37: value = 40'b1111111111111111111111111111111111111111;
						38: value = 40'b1111111111111111111111111111111111111111;
						39: value = 40'b1111111111111111111111111111111111111111;
						default: value = 40'd0;
				  endcase
				
				end
				else begin
					case(row)//black square black king
					0: value =  40'b0000000000000000000000000000000000000000;
					1: value =  40'b0000000000000000000000000000000000000000;
					2: value =  40'b0000000000000000000000000000000000000000;
					3: value =  40'b0000000000000000000000000000000000000000;
					4: value =  40'b0000000000000000000110000000000000000000;
					5: value =  40'b0000000000000000001001000000000000000000;
					6: value =  40'b0000000000000000111001110000000000000000;
					7: value =  40'b0000000000000000100000010000000000000000;
					8: value =  40'b0000000000000000111001110000000000000000;
					9: value=   40'b0000000000000000001001000000000000000000;
					10: value = 40'b0000000000000000001001000000000000000000;
					11: value = 40'b0000000000000000010000100000000000000000;
					12: value = 40'b0000000000000000100000010000000000000000;
					13: value = 40'b0000000000000001000000001000000000000000;
					14: value = 40'b0000000000000010000000000100000000000000;
					15: value = 40'b0000000000000100000000000010000000000000;
					16: value = 40'b0000000000000100000000000010000000000000;
					17: value = 40'b0000000000000010000000000100000000000000;
					18: value = 40'b0000000000000001000000001000000000000000;
					19: value = 40'b0000000000000000100000010000000000000000;
					20: value = 40'b0000000000000111110000111110000000000000;
					21: value = 40'b0000000000000100000000000010000000000000;
					22: value = 40'b0000000000000100000000000010000000000000;
					23: value = 40'b0000000000000111110000111110000000000000;
					24: value = 40'b0000000000000000010000100000000000000000;
					25: value = 40'b0000000000000000100000010000000000000000;
					26: value = 40'b0000000000000000100000010000000000000000;
					27: value = 40'b0000000000000001000000001000000000000000;
					28: value = 40'b0000000000000001000000001000000000000000;
					29: value = 40'b0000000000000010000000000100000000000000;
					30: value = 40'b0000000000000010000000000100000000000000;
					31: value = 40'b0000000000000100000000000010000000000000;
					32: value = 40'b0000000000111100000000000011110000000000;
					33: value = 40'b0000000000100000000000000000010000000000;
					34: value = 40'b0000000000100000000000000000010000000000;
					35: value = 40'b0000000000111111111111111111110000000000;
					36: value = 40'b0000000000000000000000000000000000000000;
					37: value = 40'b0000000000000000000000000000000000000000;
					38: value = 40'b0000000000000000000000000000000000000000;
					39: value = 40'b0000000000000000000000000000000000000000;
					default: value = 40'd0;
			  endcase
				end
			end
		end
		default: value = 40'd0;
	endcase
end 


endmodule 