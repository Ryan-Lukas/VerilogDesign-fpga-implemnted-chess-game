module LETTER_ROM(letteraddr,row,lettervalue);
	input [2:0] letteraddr;
	input [5:0] row;
	
	output reg [0:39] lettervalue;
	
	//all letter glyphs
	always@(*)begin
		case(letteraddr)
		3'd0: case(row) //A
			0: lettervalue =  40'b0000000000000000000000000000000000000000;
			1: lettervalue =  40'b0000000000000000000000000000000000000000;
			2: lettervalue =  40'b0000000000000000000000000000000000000000;
			3: lettervalue =  40'b0000000000000000000000000000000000000000;
			4: lettervalue =  40'b0000000000000000000000000000000000000000;
			5: lettervalue =  40'b0000000000000000000000000000000000000000;
			6: lettervalue =  40'b0000000000000000000000000000000000000000;
			7: lettervalue =  40'b0000000000000000000000000000000000000000;
			8: lettervalue =  40'b0000000000000000001111000000000000000000;
			9: lettervalue =  40'b0000000000000000011111100000000000000000;
			10: lettervalue=  40'b0000000000000000011111100000000000000000;
			11: lettervalue = 40'b0000000000000000111111110000000000000000;
			12: lettervalue = 40'b0000000000000000111111110000000000000000;
			13: lettervalue = 40'b0000000000000001111001111000000000000000;
			14: lettervalue = 40'b0000000000000001111001111000000000000000;
			15: lettervalue = 40'b0000000000000011110000111100000000000000;
			16: lettervalue = 40'b0000000000000011110000111100000000000000;
			17: lettervalue = 40'b0000000000000111110000111110000000000000;
			18: lettervalue = 40'b0000000000000111110000111110000000000000;
			19: lettervalue = 40'b0000000000001111100000011111000000000000;
			20: lettervalue = 40'b0000000000001111100000011111000000000000;
			21: lettervalue = 40'b0000000000011111000000001111100000000000;
			22: lettervalue = 40'b0000000000011111111111111111100000000000;
			23: lettervalue = 40'b0000000000111111111111111111110000000000;
			24: lettervalue = 40'b0000000000111111111111111111110000000000;
			25: lettervalue = 40'b0000000001111100000000000011111000000000;
			26: lettervalue = 40'b0000000001111100000000000011111000000000;
			27: lettervalue = 40'b0000000011111000000000000001111100000000;
			28: lettervalue = 40'b0000000011111000000000000001111100000000;
			29: lettervalue = 40'b0000000111110000000000000000111110000000;
			30: lettervalue = 40'b0000000111110000000000000000111110000000;
			31: lettervalue = 40'b0000000111110000000000000000111110000000;
			32: lettervalue = 40'b0000000000000000000000000000000000000000;
			33: lettervalue = 40'b0000000000000000000000000000000000000000;
			34: lettervalue = 40'b0000000000000000000000000000000000000000;
			35: lettervalue = 40'b0000000000000000000000000000000000000000;
			36: lettervalue = 40'b0000000000000000000000000000000000000000;
			37: lettervalue = 40'b0000000000000000000000000000000000000000;
			38: lettervalue = 40'b0000000000000000000000000000000000000000;
			39: lettervalue = 40'b0000000000000000000000000000000000000000;
			default: lettervalue = 40'd0;
		endcase 
		
		3'd1:case(row) //B
			0: lettervalue=  40'b0000000000000000000000000000000000000000;
			1: lettervalue=  40'b0000000000000000000000000000000000000000;
			2: lettervalue=  40'b0000000000000000000000000000000000000000;
			3: lettervalue=  40'b0000000000000000000000000000000000000000;
			4: lettervalue=  40'b0000000000000000000000000000000000000000;
			5: lettervalue=  40'b0000000000000000000000000000000000000000;
			6: lettervalue=  40'b0000000000000000000000000000000000000000;
			7: lettervalue=  40'b0000000000000000000000000000000000000000;
			8: lettervalue=  40'b0000000000111111111111111110000000000000;
			9: lettervalue=  40'b0000000000111111111111111111000000000000;
			10:lettervalue=  40'b0000000000111111111111111111100000000000;
			11:lettervalue = 40'b0000000000111100000000001111110000000000;
			12:lettervalue = 40'b0000000000111100000000000111111000000000;
			13:lettervalue = 40'b0000000000111100000000000011111000000000;
			14:lettervalue = 40'b0000000000111100000000000011111000000000;
			15:lettervalue = 40'b0000000000111100000000000011111000000000;
			16:lettervalue = 40'b0000000000111100000000000011111000000000;
			17:lettervalue = 40'b0000000000111100000000000111110000000000;
			18:lettervalue = 40'b0000000000111100000000001111100000000000;
			19:lettervalue = 40'b0000000000111111111111111111000000000000;
			20:lettervalue = 40'b0000000000111111111111111111000000000000;
			21:lettervalue = 40'b0000000000111100000000001111100000000000;
			22:lettervalue = 40'b0000000000111100000000000111110000000000;
			23:lettervalue = 40'b0000000000111100000000000011111000000000;
			24:lettervalue = 40'b0000000000111100000000000001111000000000;
			25:lettervalue = 40'b0000000000111100000000000001111000000000;
			26:lettervalue = 40'b0000000000111100000000000001111000000000;
			27:lettervalue = 40'b0000000000111100000000000001111000000000;
			28:lettervalue = 40'b0000000000111100000000000011111000000000;
			29:lettervalue = 40'b0000000000111111111111111111110000000000;
			30:lettervalue = 40'b0000000000111111111111111111100000000000;
			31:lettervalue = 40'b0000000000111111111111111111000000000000;
			32:lettervalue = 40'b0000000000000000000000000000000000000000;
			33:lettervalue = 40'b0000000000000000000000000000000000000000;
			34:lettervalue = 40'b0000000000000000000000000000000000000000;
			35:lettervalue = 40'b0000000000000000000000000000000000000000;
			36:lettervalue = 40'b0000000000000000000000000000000000000000;
			37:lettervalue = 40'b0000000000000000000000000000000000000000;
			38:lettervalue = 40'b0000000000000000000000000000000000000000;
			39:lettervalue = 40'b0000000000000000000000000000000000000000;
			default: lettervalue = 40'd0;
		endcase 
		
		3'd2:case(row) //C
			0: lettervalue =  40'b0000000000000000000000000000000000000000;
			1: lettervalue =  40'b0000000000000000000000000000000000000000;
			2: lettervalue =  40'b0000000000000000000000000000000000000000;
			3: lettervalue =  40'b0000000000000000000000000000000000000000;
			4: lettervalue =  40'b0000000000000000000000000000000000000000;
			5: lettervalue =  40'b0000000000000000000000000000000000000000;
			6: lettervalue =  40'b0000000000000000000000000000000000000000;
			7: lettervalue =  40'b0000000000000000000000000000000000000000;
			8: lettervalue =  40'b0000000000111111111111111111110000000000;
			9: lettervalue =  40'b0000000000111111111111111111110000000000;
			10: lettervalue=  40'b0000000000111111111111111111110000000000;
			11: lettervalue = 40'b0000000000111110000000000011110000000000;
			12: lettervalue = 40'b0000000000111110000000000011110000000000;
			13: lettervalue = 40'b0000000000111110000000000011110000000000;
			14: lettervalue = 40'b0000000000111110000000000011110000000000;
			15: lettervalue = 40'b0000000000111110000000000000000000000000;
			16: lettervalue = 40'b0000000000111110000000000000000000000000;
			17: lettervalue = 40'b0000000000111110000000000000000000000000;
			18: lettervalue = 40'b0000000000111110000000000000000000000000;
			19: lettervalue = 40'b0000000000111110000000000000000000000000;
			20: lettervalue = 40'b0000000000111110000000000000000000000000;
			21: lettervalue = 40'b0000000000111110000000000000000000000000;
			22: lettervalue = 40'b0000000000111110000000000000000000000000;
			23: lettervalue = 40'b0000000000111110000000000000000000000000;
			24: lettervalue = 40'b0000000000111110000000000000000000000000;
			25: lettervalue = 40'b0000000000111110000000000011110000000000;
			26: lettervalue = 40'b0000000000111110000000000011110000000000;
			27: lettervalue = 40'b0000000000111110000000000011110000000000;
			28: lettervalue = 40'b0000000000111110000000000011110000000000;
			29: lettervalue = 40'b0000000000111111111111111111110000000000;
			30: lettervalue = 40'b0000000000111111111111111111110000000000;
			31: lettervalue = 40'b0000000000111111111111111111110000000000;
			32: lettervalue = 40'b0000000000000000000000000000000000000000;
			33: lettervalue = 40'b0000000000000000000000000000000000000000;
			34: lettervalue = 40'b0000000000000000000000000000000000000000;
			35: lettervalue = 40'b0000000000000000000000000000000000000000;
			36: lettervalue = 40'b0000000000000000000000000000000000000000;
			37: lettervalue = 40'b0000000000000000000000000000000000000000;
			38: lettervalue = 40'b0000000000000000000000000000000000000000;
			39: lettervalue = 40'b0000000000000000000000000000000000000000;
			default: lettervalue = 40'd0;
		endcase 
		
		3'd3:case(row) //D
			0: lettervalue =  40'b0000000000000000000000000000000000000000;
			1: lettervalue =  40'b0000000000000000000000000000000000000000;
			2: lettervalue =  40'b0000000000000000000000000000000000000000;
			3: lettervalue =  40'b0000000000000000000000000000000000000000;
			4: lettervalue =  40'b0000000000000000000000000000000000000000;
			5: lettervalue =  40'b0000000000000000000000000000000000000000;
			6: lettervalue =  40'b0000000000000000000000000000000000000000;
			7: lettervalue =  40'b0000000000000000000000000000000000000000;
			8: lettervalue =  40'b0000000000111111111111100000000000000000;
			9: lettervalue =  40'b0000000000111111111111110000000000000000;
			10: lettervalue=  40'b0000000000111111111111111000000000000000;
			11: lettervalue = 40'b0000000000111111111111111100000000000000;
			12: lettervalue = 40'b0000000000111100000000011110000000000000;
			13: lettervalue = 40'b0000000000111100000000001111000000000000;
			14: lettervalue = 40'b0000000000111100000000000111100000000000;
			15: lettervalue = 40'b0000000000111100000000000111100000000000;
			16: lettervalue = 40'b0000000000111100000000000111100000000000;
			17: lettervalue = 40'b0000000000111100000000000111100000000000;
			18: lettervalue = 40'b0000000000111100000000000111100000000000;
			19: lettervalue = 40'b0000000000111100000000000111100000000000;
			20: lettervalue = 40'b0000000000111100000000000111100000000000;
			21: lettervalue = 40'b0000000000111100000000000111100000000000;
			22: lettervalue = 40'b0000000000111100000000000111100000000000;
			23: lettervalue = 40'b0000000000111100000000000111100000000000;
			24: lettervalue = 40'b0000000000111100000000000111100000000000;
			25: lettervalue = 40'b0000000000111100000000000111100000000000;
			26: lettervalue = 40'b0000000000111100000000001111000000000000;
			27: lettervalue = 40'b0000000000111100000000011110000000000000;
			28: lettervalue = 40'b0000000000111111111111111100000000000000;
			29: lettervalue = 40'b0000000000111111111111111000000000000000;
			30: lettervalue = 40'b0000000000111111111111110000000000000000;
			31: lettervalue = 40'b0000000000111111111111100000000000000000;
			32: lettervalue = 40'b0000000000000000000000000000000000000000;
			33: lettervalue = 40'b0000000000000000000000000000000000000000;
			34: lettervalue = 40'b0000000000000000000000000000000000000000;
			35: lettervalue = 40'b0000000000000000000000000000000000000000;
			36: lettervalue = 40'b0000000000000000000000000000000000000000;
			37: lettervalue = 40'b0000000000000000000000000000000000000000;
			38: lettervalue = 40'b0000000000000000000000000000000000000000;
			39: lettervalue = 40'b0000000000000000000000000000000000000000;
			default: lettervalue = 40'd0;
		endcase 
		
		3'd4:case(row) //E
			0: lettervalue =  40'b0000000000000000000000000000000000000000;
			1: lettervalue =  40'b0000000000000000000000000000000000000000;
			2: lettervalue =  40'b0000000000000000000000000000000000000000;
			3: lettervalue =  40'b0000000000000000000000000000000000000000;
			4: lettervalue =  40'b0000000000000000000000000000000000000000;
			5: lettervalue =  40'b0000000000000000000000000000000000000000;
			6: lettervalue =  40'b0000000000000000000000000000000000000000;
			7: lettervalue =  40'b0000000000000000000000000000000000000000;
			8: lettervalue =  40'b0000000000111111111111111111100000000000;
			9: lettervalue =  40'b0000000000111111111111111111100000000000;
			10: lettervalue=  40'b0000000000111111111111111111100000000000;
			11: lettervalue = 40'b0000000000111110000000000000000000000000;
			12: lettervalue = 40'b0000000000111110000000000000000000000000;
			13: lettervalue = 40'b0000000000111110000000000000000000000000;
			14: lettervalue = 40'b0000000000111110000000000000000000000000;
			15: lettervalue = 40'b0000000000111110000000000000000000000000;
			16: lettervalue = 40'b0000000000111110000000000000000000000000;
			17: lettervalue = 40'b0000000000111110000000000000000000000000;
			18: lettervalue = 40'b0000000000111111111111111110000000000000;
			19: lettervalue = 40'b0000000000111111111111111110000000000000;
			20: lettervalue = 40'b0000000000111111111111111110000000000000;
			21: lettervalue = 40'b0000000000111110000000000000000000000000;
			22: lettervalue = 40'b0000000000111110000000000000000000000000;
			23: lettervalue = 40'b0000000000111110000000000000000000000000;
			24: lettervalue = 40'b0000000000111110000000000000000000000000;
			25: lettervalue = 40'b0000000000111110000000000000000000000000;
			26: lettervalue = 40'b0000000000111110000000000000000000000000;
			27: lettervalue = 40'b0000000000111110000000000000000000000000;
			28: lettervalue = 40'b0000000000111110000000000000000000000000;
			29: lettervalue = 40'b0000000000111111111111111111100000000000;
			30: lettervalue = 40'b0000000000111111111111111111100000000000;
			31: lettervalue = 40'b0000000000111111111111111111100000000000;
			32: lettervalue = 40'b0000000000000000000000000000000000000000;
			33: lettervalue = 40'b0000000000000000000000000000000000000000;
			34: lettervalue = 40'b0000000000000000000000000000000000000000;
			35: lettervalue = 40'b0000000000000000000000000000000000000000;
			36: lettervalue = 40'b0000000000000000000000000000000000000000;
			37: lettervalue = 40'b0000000000000000000000000000000000000000;
			38: lettervalue = 40'b0000000000000000000000000000000000000000;
			39: lettervalue = 40'b0000000000000000000000000000000000000000;
			default: lettervalue = 40'd0;
		endcase 
		
		3'd5:case(row) //F
			0: lettervalue =  40'b0000000000000000000000000000000000000000;
			1: lettervalue =  40'b0000000000000000000000000000000000000000;
			2: lettervalue =  40'b0000000000000000000000000000000000000000;
			3: lettervalue =  40'b0000000000000000000000000000000000000000;
			4: lettervalue =  40'b0000000000000000000000000000000000000000;
			5: lettervalue =  40'b0000000000000000000000000000000000000000;
			6: lettervalue =  40'b0000000000000000000000000000000000000000;
			7: lettervalue =  40'b0000000000000000000000000000000000000000;
			8: lettervalue =  40'b0000000000011111111111111110000000000000;
			9: lettervalue =  40'b0000000000011111111111111110000000000000;
			10: lettervalue=  40'b0000000000011111111111111110000000000000;
			11: lettervalue = 40'b0000000000011111000000000000000000000000;
			12: lettervalue = 40'b0000000000011111000000000000000000000000;
			13: lettervalue = 40'b0000000000011111000000000000000000000000;
			14: lettervalue = 40'b0000000000011111000000000000000000000000;
			15: lettervalue = 40'b0000000000011111000000000000000000000000;
			16: lettervalue = 40'b0000000000011111000000000000000000000000;
			17: lettervalue = 40'b0000000000011111111111111000000000000000;
			18: lettervalue = 40'b0000000000011111111111111000000000000000;
			19: lettervalue = 40'b0000000000011111111111111000000000000000;
			20: lettervalue = 40'b0000000000011111000000000000000000000000;
			21: lettervalue = 40'b0000000000011111000000000000000000000000;
			22: lettervalue = 40'b0000000000011111000000000000000000000000;
			23: lettervalue = 40'b0000000000011111000000000000000000000000;
			24: lettervalue = 40'b0000000000011111000000000000000000000000;
			25: lettervalue = 40'b0000000000011111000000000000000000000000;
			26: lettervalue = 40'b0000000000011111000000000000000000000000;
			27: lettervalue = 40'b0000000000011111000000000000000000000000;
			28: lettervalue = 40'b0000000000011111000000000000000000000000;
			29: lettervalue = 40'b0000000000011111000000000000000000000000;
			30: lettervalue = 40'b0000000000011111000000000000000000000000;
			31: lettervalue = 40'b0000000000011111000000000000000000000000;
			32: lettervalue = 40'b0000000000000000000000000000000000000000;
			33: lettervalue = 40'b0000000000000000000000000000000000000000;
			34: lettervalue = 40'b0000000000000000000000000000000000000000;
			35: lettervalue = 40'b0000000000000000000000000000000000000000;
			36: lettervalue = 40'b0000000000000000000000000000000000000000;
			37: lettervalue = 40'b0000000000000000000000000000000000000000;
			38: lettervalue = 40'b0000000000000000000000000000000000000000;
			39: lettervalue = 40'b0000000000000000000000000000000000000000;
			default: lettervalue = 40'd0;
		endcase 
		
		3'd6:case(row) //G
			0: lettervalue =  40'b0000000000000000000000000000000000000000;
			1: lettervalue =  40'b0000000000000000000000000000000000000000;
			2: lettervalue =  40'b0000000000000000000000000000000000000000;
			3: lettervalue =  40'b0000000000000000000000000000000000000000;
			4: lettervalue =  40'b0000000000000000000000000000000000000000;
			5: lettervalue =  40'b0000000000000000000000000000000000000000;
			6: lettervalue =  40'b0000000000000000000000000000000000000000;
			7: lettervalue =  40'b0000000000000000000000000000000000000000;
			8: lettervalue =  40'b0000000000111111111111111111110000000000;
			9: lettervalue =  40'b0000000000111111111111111111110000000000;
			10: lettervalue=  40'b0000000000111111111111111111110000000000;
			11: lettervalue = 40'b0000000000111110000000000011110000000000;
			12: lettervalue = 40'b0000000000111110000000000011110000000000;
			13: lettervalue = 40'b0000000000111110000000000011110000000000;
			14: lettervalue = 40'b0000000000111110000000000011110000000000;
			15: lettervalue = 40'b0000000000111110000000000000000000000000;
			16: lettervalue = 40'b0000000000111110000000000000000000000000;
			17: lettervalue = 40'b0000000000111110000000000000000000000000;
			18: lettervalue = 40'b0000000000111110000000000000000000000000;
			19: lettervalue = 40'b0000000000111110000011111111110000000000;
			20: lettervalue = 40'b0000000000111110000011111111110000000000;
			21: lettervalue = 40'b0000000000111110000011111111110000000000;
			22: lettervalue = 40'b0000000000111110000000000011110000000000;
			23: lettervalue = 40'b0000000000111110000000000011110000000000;
			24: lettervalue = 40'b0000000000111110000000000011110000000000;
			25: lettervalue = 40'b0000000000111110000000000011110000000000;
			26: lettervalue = 40'b0000000000111110000000000011110000000000;
			27: lettervalue = 40'b0000000000111110000000000011110000000000;
			28: lettervalue = 40'b0000000000111110000000000011110000000000;
			29: lettervalue = 40'b0000000000111111111111111111110000000000;
			30: lettervalue = 40'b0000000000111111111111111111110000000000;
			31: lettervalue = 40'b0000000000111111111111111111110000000000;
			32: lettervalue = 40'b0000000000000000000000000000000000000000;
			33: lettervalue = 40'b0000000000000000000000000000000000000000;
			34: lettervalue = 40'b0000000000000000000000000000000000000000;
			35: lettervalue = 40'b0000000000000000000000000000000000000000;
			36: lettervalue = 40'b0000000000000000000000000000000000000000;
			37: lettervalue = 40'b0000000000000000000000000000000000000000;
			38: lettervalue = 40'b0000000000000000000000000000000000000000;
			39: lettervalue = 40'b0000000000000000000000000000000000000000;
			default: lettervalue = 40'd0;
		endcase 
		
		3'd7:case(row) //H
			0: lettervalue =  40'b0000000000000000000000000000000000000000;
			1: lettervalue =  40'b0000000000000000000000000000000000000000;
			2: lettervalue =  40'b0000000000000000000000000000000000000000;
			3: lettervalue =  40'b0000000000000000000000000000000000000000;
			4: lettervalue =  40'b0000000000000000000000000000000000000000;
			5: lettervalue =  40'b0000000000000000000000000000000000000000;
			6: lettervalue =  40'b0000000000000000000000000000000000000000;
			7: lettervalue =  40'b0000000000000000000000000000000000000000;
			8: lettervalue =  40'b0000000000011111000000001111100000000000;
			9: lettervalue =  40'b0000000000011111000000001111100000000000;
			10: lettervalue=  40'b0000000000011111000000001111100000000000;
			11: lettervalue = 40'b0000000000011111000000001111100000000000;
			12: lettervalue = 40'b0000000000011111000000001111100000000000;
			13: lettervalue = 40'b0000000000011111000000001111100000000000;
			14: lettervalue = 40'b0000000000011111000000001111100000000000;
			15: lettervalue = 40'b0000000000011111000000001111100000000000;
			16: lettervalue = 40'b0000000000011111000000001111100000000000;
			17: lettervalue = 40'b0000000000011111111111111111100000000000;
			18: lettervalue = 40'b0000000000011111111111111111100000000000;
			19: lettervalue = 40'b0000000000011111111111111111100000000000;
			20: lettervalue = 40'b0000000000011111111111111111100000000000;
			21: lettervalue = 40'b0000000000011111000000001111100000000000;
			22: lettervalue = 40'b0000000000011111000000001111100000000000;
			23: lettervalue = 40'b0000000000011111000000001111100000000000;
			24: lettervalue = 40'b0000000000011111000000001111100000000000;
			25: lettervalue = 40'b0000000000011111000000001111100000000000;
			26: lettervalue = 40'b0000000000011111000000001111100000000000;
			27: lettervalue = 40'b0000000000011111000000001111100000000000;
			28: lettervalue = 40'b0000000000011111000000001111100000000000;
			29: lettervalue = 40'b0000000000011111000000001111100000000000;
			30: lettervalue = 40'b0000000000011111000000001111100000000000;
			31: lettervalue = 40'b0000000000011111000000001111100000000000;
			32: lettervalue = 40'b0000000000000000000000000000000000000000;
			33: lettervalue = 40'b0000000000000000000000000000000000000000;
			34: lettervalue = 40'b0000000000000000000000000000000000000000;
			35: lettervalue = 40'b0000000000000000000000000000000000000000;
			36: lettervalue = 40'b0000000000000000000000000000000000000000;
			37: lettervalue = 40'b0000000000000000000000000000000000000000;
			38: lettervalue = 40'b0000000000000000000000000000000000000000;
			39: lettervalue = 40'b0000000000000000000000000000000000000000;
			default: lettervalue = 40'd0;
		endcase 
		
		
		default: lettervalue = 40'd0;
		
		endcase
	end

endmodule
