module NUMBER_ROM(numberaddr,row,numbervalue);
input [2:0] numberaddr;
input [5:0] row;
output reg [0:39] numbervalue;


always@(*)begin
	//number glyph selection
	case(numberaddr)
		3'd0:case(row) //8
			0: numbervalue =  40'b0000000000000000000000000000000000000000;
			1: numbervalue =  40'b0000000000000000000000000000000000000000;
			2: numbervalue =  40'b0000000000000000000000000000000000000000;
			3: numbervalue =  40'b0000000000000000000000000000000000000000;
			4: numbervalue =  40'b0000000000000000000000000000000000000000;
			5: numbervalue =  40'b0000000000000000000000000000000000000000;
			6: numbervalue =  40'b0000000000000000000000000000000000000000;
			7: numbervalue =  40'b0000000000000000000000000000000000000000;
			8: numbervalue =  40'b0000000000111111111111111111000000000000;
			9: numbervalue =  40'b0000000000111111111111111111000000000000;
			10: numbervalue=  40'b0000000000111111111111111111000000000000;
			11: numbervalue = 40'b0000000000111110000000011111000000000000;
			12: numbervalue = 40'b0000000000111110000000011111000000000000;
			13: numbervalue = 40'b0000000000111110000000011111000000000000;
			14: numbervalue = 40'b0000000000111110000000011111000000000000;
			15: numbervalue = 40'b0000000000111110000000011111000000000000;
			16: numbervalue = 40'b0000000000111110000000011111000000000000;
			17: numbervalue = 40'b0000000000111110000000011111000000000000;
			18: numbervalue = 40'b0000000000111111111111111111000000000000;
			19: numbervalue = 40'b0000000000111111111111111111000000000000;
			20: numbervalue = 40'b0000000000111111111111111111000000000000;
			21: numbervalue = 40'b0000000000111110000000011111000000000000;
			22: numbervalue = 40'b0000000000111110000000011111000000000000;
			23: numbervalue = 40'b0000000000111110000000011111000000000000;
			24: numbervalue = 40'b0000000000111110000000011111000000000000;
			25: numbervalue = 40'b0000000000111110000000011111000000000000;
			26: numbervalue = 40'b0000000000111110000000011111000000000000;
			27: numbervalue = 40'b0000000000111110000000011111000000000000;
			28: numbervalue = 40'b0000000000111110000000011111000000000000;
			29: numbervalue = 40'b0000000000111111111111111111000000000000;
			30: numbervalue = 40'b0000000000111111111111111111000000000000;
			31: numbervalue = 40'b0000000000111111111111111111000000000000;
			32: numbervalue = 40'b0000000000000000000000000000000000000000;
			33: numbervalue = 40'b0000000000000000000000000000000000000000;
			34: numbervalue = 40'b0000000000000000000000000000000000000000;
			35: numbervalue = 40'b0000000000000000000000000000000000000000;
			36: numbervalue = 40'b0000000000000000000000000000000000000000;
			37: numbervalue = 40'b0000000000000000000000000000000000000000;
			38: numbervalue = 40'b0000000000000000000000000000000000000000;
			39: numbervalue = 40'b0000000000000000000000000000000000000000;
			default: numbervalue = 40'd0;
		endcase 
		
			3'd1:case(row) //7
			0: numbervalue =  40'b0000000000000000000000000000000000000000;
			1: numbervalue =  40'b0000000000000000000000000000000000000000;
			2: numbervalue =  40'b0000000000000000000000000000000000000000;
			3: numbervalue =  40'b0000000000000000000000000000000000000000;
			4: numbervalue =  40'b0000000000000000000000000000000000000000;
			5: numbervalue =  40'b0000000000000000000000000000000000000000;
			6: numbervalue =  40'b0000000000000000000000000000000000000000;
			7: numbervalue =  40'b0000000000000000000000000000000000000000;
			8: numbervalue =  40'b0000000000011111111111111111100000000000;
			9: numbervalue =  40'b0000000000011111111111111111100000000000;
			10: numbervalue=  40'b0000000000011111111111111111100000000000;
			11: numbervalue = 40'b0000000000000000000000001111100000000000;
			12: numbervalue = 40'b0000000000000000000000001111100000000000;
			13: numbervalue = 40'b0000000000000000000000001111100000000000;
			14: numbervalue = 40'b0000000000000000000000011111000000000000;
			15: numbervalue = 40'b0000000000000000000000011111000000000000;
			16: numbervalue = 40'b0000000000000000000000111110000000000000;
			17: numbervalue = 40'b0000000000000000000000111110000000000000;
			18: numbervalue = 40'b0000000000000000000001111100000000000000;
			19: numbervalue = 40'b0000000000000000000001111100000000000000;
			20: numbervalue = 40'b0000000000000000000011111000000000000000;
			21: numbervalue = 40'b0000000000000000000011111000000000000000;
			22: numbervalue = 40'b0000000000000000000111110000000000000000;
			23: numbervalue = 40'b0000000000000000000111110000000000000000;
			24: numbervalue = 40'b0000000000000000001111100000000000000000;
			25: numbervalue = 40'b0000000000000000001111100000000000000000;
			26: numbervalue = 40'b0000000000000000011111000000000000000000;
			27: numbervalue = 40'b0000000000000000011111000000000000000000;
			28: numbervalue = 40'b0000000000000000111110000000000000000000;
			29: numbervalue = 40'b0000000000000000111110000000000000000000;
			30: numbervalue = 40'b0000000000000001111100000000000000000000;
			31: numbervalue = 40'b0000000000000001111100000000000000000000;
			32: numbervalue = 40'b0000000000000000000000000000000000000000;
			33: numbervalue = 40'b0000000000000000000000000000000000000000;
			34: numbervalue = 40'b0000000000000000000000000000000000000000;
			35: numbervalue = 40'b0000000000000000000000000000000000000000;
			36: numbervalue = 40'b0000000000000000000000000000000000000000;
			37: numbervalue = 40'b0000000000000000000000000000000000000000;
			38: numbervalue = 40'b0000000000000000000000000000000000000000;
			39: numbervalue = 40'b0000000000000000000000000000000000000000;
			default: numbervalue = 40'd0;
		endcase
		
		3'd2:case(row) //6
			0: numbervalue =  40'b0000000000000000000000000000000000000000;
			1: numbervalue =  40'b0000000000000000000000000000000000000000;
			2: numbervalue =  40'b0000000000000000000000000000000000000000;
			3: numbervalue =  40'b0000000000000000000000000000000000000000;
			4: numbervalue =  40'b0000000000000000000000000000000000000000;
			5: numbervalue =  40'b0000000000000000000000000000000000000000;
			6: numbervalue =  40'b0000000000000000000000000000000000000000;
			7: numbervalue =  40'b0000000000000000000000000000000000000000;
			8: numbervalue =  40'b0000000000011111111111111111100000000000;
			9: numbervalue =  40'b0000000000011111111111111111100000000000;
			10: numbervalue=  40'b0000000000011111111111111111100000000000;
			11: numbervalue = 40'b0000000000011110000000000000000000000000;
			12: numbervalue = 40'b0000000000011110000000000000000000000000;
			13: numbervalue = 40'b0000000000011110000000000000000000000000;
			14: numbervalue = 40'b0000000000011110000000000000000000000000;
			15: numbervalue = 40'b0000000000011110000000000000000000000000;
			16: numbervalue = 40'b0000000000011110000000000000000000000000;
			17: numbervalue = 40'b0000000000011110000000000000000000000000;
			18: numbervalue = 40'b0000000000011111111111111111100000000000;
			19: numbervalue = 40'b0000000000011111111111111111100000000000;
			20: numbervalue = 40'b0000000000011111111111111111100000000000;
			21: numbervalue = 40'b0000000000011110000000000111100000000000;
			22: numbervalue = 40'b0000000000011110000000000111100000000000;
			23: numbervalue = 40'b0000000000011110000000000111100000000000;
			24: numbervalue = 40'b0000000000011110000000000111100000000000;
			25: numbervalue = 40'b0000000000011110000000000111100000000000;
			26: numbervalue = 40'b0000000000011110000000000111100000000000;
			27: numbervalue = 40'b0000000000011110000000000111100000000000;
			28: numbervalue = 40'b0000000000011110000000000111100000000000;
			29: numbervalue = 40'b0000000000011111111111111111100000000000;
			30: numbervalue = 40'b0000000000011111111111111111100000000000;
			31: numbervalue = 40'b0000000000011111111111111111100000000000;
			32: numbervalue = 40'b0000000000000000000000000000000000000000;
			33: numbervalue = 40'b0000000000000000000000000000000000000000;
			34: numbervalue = 40'b0000000000000000000000000000000000000000;
			35: numbervalue = 40'b0000000000000000000000000000000000000000;
			36: numbervalue = 40'b0000000000000000000000000000000000000000;
			37: numbervalue = 40'b0000000000000000000000000000000000000000;
			38: numbervalue = 40'b0000000000000000000000000000000000000000;
			39: numbervalue = 40'b0000000000000000000000000000000000000000;
			default: numbervalue = 40'd0;
		endcase 
		
		3'd3:case(row) //5
			0: numbervalue =  40'b0000000000000000000000000000000000000000;
			1: numbervalue =  40'b0000000000000000000000000000000000000000;
			2: numbervalue =  40'b0000000000000000000000000000000000000000;
			3: numbervalue =  40'b0000000000000000000000000000000000000000;
			4: numbervalue =  40'b0000000000000000000000000000000000000000;
			5: numbervalue =  40'b0000000000000000000000000000000000000000;
			6: numbervalue =  40'b0000000000000000000000000000000000000000;
			7: numbervalue =  40'b0000000000000000000000000000000000000000;
			8: numbervalue =  40'b0000000000011111111111111111100000000000;
			9: numbervalue =  40'b0000000000011111111111111111100000000000;
			10: numbervalue=  40'b0000000000011111111111111111100000000000;
			11: numbervalue = 40'b0000000000011110000000000000000000000000;
			12: numbervalue = 40'b0000000000011110000000000000000000000000;
			13: numbervalue = 40'b0000000000011110000000000000000000000000;
			14: numbervalue = 40'b0000000000011110000000000000000000000000;
			15: numbervalue = 40'b0000000000011110000000000000000000000000;
			16: numbervalue = 40'b0000000000011110000000000000000000000000;
			17: numbervalue = 40'b0000000000011110000000000000000000000000;
			18: numbervalue = 40'b0000000000011110000000000000000000000000;
			19: numbervalue = 40'b0000000000011111111111111111100000000000;
			20: numbervalue = 40'b0000000000011111111111111111100000000000;
			21: numbervalue = 40'b0000000000011111111111111111100000000000;
			22: numbervalue = 40'b0000000000000000000000000111100000000000;
			23: numbervalue = 40'b0000000000000000000000000111100000000000;
			24: numbervalue = 40'b0000000000000000000000000111100000000000;
			25: numbervalue = 40'b0000000000000000000000000111100000000000;
			26: numbervalue = 40'b0000000000000000000000000111100000000000;
			27: numbervalue = 40'b0000000000000000000000000111100000000000;
			28: numbervalue = 40'b0000000000000000000000000111100000000000;
			29: numbervalue = 40'b0000000000011111111111111111100000000000;
			30: numbervalue = 40'b0000000000011111111111111111100000000000;
			31: numbervalue = 40'b0000000000011111111111111111100000000000;
			32: numbervalue = 40'b0000000000000000000000000000000000000000;
			33: numbervalue = 40'b0000000000000000000000000000000000000000;
			34: numbervalue = 40'b0000000000000000000000000000000000000000;
			35: numbervalue = 40'b0000000000000000000000000000000000000000;
			36: numbervalue = 40'b0000000000000000000000000000000000000000;
			37: numbervalue = 40'b0000000000000000000000000000000000000000;
			38: numbervalue = 40'b0000000000000000000000000000000000000000;
			39: numbervalue = 40'b0000000000000000000000000000000000000000;
			default: numbervalue = 40'd0;
		endcase
		
		3'd4: case(row) //4
			0: numbervalue =  40'b0000000000000000000000000000000000000000;
			1: numbervalue =  40'b0000000000000000000000000000000000000000;
			2: numbervalue =  40'b0000000000000000000000000000000000000000;
			3: numbervalue =  40'b0000000000000000000000000000000000000000;
			4: numbervalue =  40'b0000000000000000000000000000000000000000;
			5: numbervalue =  40'b0000000000000000000000000000000000000000;
			6: numbervalue =  40'b0000000000000000000000000000000000000000;
			7: numbervalue =  40'b0000000000000000000000000000000000000000;
			8: numbervalue =  40'b0000000000011111000001111100000000000000;
			9: numbervalue =  40'b0000000000011111000001111100000000000000;
			10: numbervalue=  40'b0000000000011111000001111100000000000000;
			11: numbervalue = 40'b0000000000011111000001111100000000000000;
			12: numbervalue = 40'b0000000000011111000001111100000000000000;
			13: numbervalue = 40'b0000000000011111000001111100000000000000;
			14: numbervalue = 40'b0000000000011111000001111100000000000000;
			15: numbervalue = 40'b0000000000011111000001111100000000000000;
			16: numbervalue = 40'b0000000000011111000001111100000000000000;
			17: numbervalue = 40'b0000000000011111000001111100000000000000;
			18: numbervalue = 40'b0000000000011111000001111100000000000000;
			19: numbervalue = 40'b0000000000011111000001111100000000000000;
			20: numbervalue = 40'b0000000000011111000001111100000000000000;
			21: numbervalue = 40'b0000000000011111111111111111100000000000;
			22: numbervalue = 40'b0000000000011111111111111111100000000000;
			23: numbervalue = 40'b0000000000011111111111111111100000000000;
			24: numbervalue = 40'b0000000000000000000001111100000000000000;
			25: numbervalue = 40'b0000000000000000000001111100000000000000;
			26: numbervalue = 40'b0000000000000000000001111100000000000000;
			27: numbervalue = 40'b0000000000000000000001111100000000000000;
			28: numbervalue = 40'b0000000000000000000001111100000000000000;
			29: numbervalue = 40'b0000000000000000000001111100000000000000;
			30: numbervalue = 40'b0000000000000000000001111100000000000000;
			31: numbervalue = 40'b0000000000000000000001111100000000000000;
			32: numbervalue = 40'b0000000000000000000000000000000000000000;
			33: numbervalue = 40'b0000000000000000000000000000000000000000;
			34: numbervalue = 40'b0000000000000000000000000000000000000000;
			35: numbervalue = 40'b0000000000000000000000000000000000000000;
			36: numbervalue = 40'b0000000000000000000000000000000000000000;
			37: numbervalue = 40'b0000000000000000000000000000000000000000;
			38: numbervalue = 40'b0000000000000000000000000000000000000000;
			39: numbervalue = 40'b0000000000000000000000000000000000000000;
			default: numbervalue = 40'd0;
		endcase
		
			3'd5:case(row) //3
			0: numbervalue =  40'b0000000000000000000000000000000000000000;
			1: numbervalue =  40'b0000000000000000000000000000000000000000;
			2: numbervalue =  40'b0000000000000000000000000000000000000000;
			3: numbervalue =  40'b0000000000000000000000000000000000000000;
			4: numbervalue =  40'b0000000000000000000000000000000000000000;
			5: numbervalue =  40'b0000000000000000000000000000000000000000;
			6: numbervalue =  40'b0000000000000000000000000000000000000000;
			7: numbervalue =  40'b0000000000000000000000000000000000000000;
			8: numbervalue =  40'b0000000000011111111111111111100000000000;
			9: numbervalue =  40'b0000000000011111111111111111100000000000;
			10: numbervalue=  40'b0000000000011111111111111111100000000000;
			11: numbervalue = 40'b0000000000000000000000001111100000000000;
			12: numbervalue = 40'b0000000000000000000000001111100000000000;
			13: numbervalue = 40'b0000000000000000000000001111100000000000;
			14: numbervalue = 40'b0000000000000000000000001111100000000000;
			15: numbervalue = 40'b0000000000000000000000001111100000000000;
			16: numbervalue = 40'b0000000000000000000000001111100000000000;
			17: numbervalue = 40'b0000000000000000000000001111100000000000;
			18: numbervalue = 40'b0000000000000000000000001111100000000000;
			19: numbervalue = 40'b0000000000011111111111111111100000000000;
			20: numbervalue = 40'b0000000000011111111111111111100000000000;
			21: numbervalue = 40'b0000000000011111111111111111100000000000;
			22: numbervalue = 40'b0000000000000000000000001111100000000000;
			23: numbervalue = 40'b0000000000000000000000001111100000000000;
			24: numbervalue = 40'b0000000000000000000000001111100000000000;
			25: numbervalue = 40'b0000000000000000000000001111100000000000;
			26: numbervalue = 40'b0000000000000000000000001111100000000000;
			27: numbervalue = 40'b0000000000000000000000001111100000000000;
			28: numbervalue = 40'b0000000000000000000000001111100000000000;
			29: numbervalue = 40'b0000000000011111111111111111100000000000;
			30: numbervalue = 40'b0000000000011111111111111111100000000000;
			31: numbervalue = 40'b0000000000011111111111111111100000000000;
			32: numbervalue = 40'b0000000000000000000000000000000000000000;
			33: numbervalue = 40'b0000000000000000000000000000000000000000;
			34: numbervalue = 40'b0000000000000000000000000000000000000000;
			35: numbervalue = 40'b0000000000000000000000000000000000000000;
			36: numbervalue = 40'b0000000000000000000000000000000000000000;
			37: numbervalue = 40'b0000000000000000000000000000000000000000;
			38: numbervalue = 40'b0000000000000000000000000000000000000000;
			39: numbervalue = 40'b0000000000000000000000000000000000000000;
			default: numbervalue = 40'd0;
		endcase 
		
		3'd6:case(row) //2
			0: numbervalue =  40'b0000000000000000000000000000000000000000;
			1: numbervalue =  40'b0000000000000000000000000000000000000000;
			2: numbervalue =  40'b0000000000000000000000000000000000000000;
			3: numbervalue =  40'b0000000000000000000000000000000000000000;
			4: numbervalue =  40'b0000000000000000000000000000000000000000;
			5: numbervalue =  40'b0000000000000000000000000000000000000000;
			6: numbervalue =  40'b0000000000000000000000000000000000000000;
			7: numbervalue =  40'b0000000000000000000000000000000000000000;
			8: numbervalue =  40'b0000000000111111111111111111000000000000;
			9: numbervalue =  40'b0000000000111111111111111111000000000000;
			10: numbervalue=  40'b0000000000111111111111111111000000000000;
			11: numbervalue = 40'b0000000000000000000000001111000000000000;
			12: numbervalue = 40'b0000000000000000000000001111000000000000;
			13: numbervalue = 40'b0000000000000000000000001111000000000000;
			14: numbervalue = 40'b0000000000000000000000001111000000000000;
			15: numbervalue = 40'b0000000000000000000000001111000000000000;
			16: numbervalue = 40'b0000000000000000000000001111000000000000;
			17: numbervalue = 40'b0000000000000000000000001111000000000000;
			18: numbervalue = 40'b0000000000111111111111111111000000000000;
			19: numbervalue = 40'b0000000000111111111111111111000000000000;
			20: numbervalue = 40'b0000000000111111111111111111000000000000;
			21: numbervalue = 40'b0000000000111100000000000000000000000000;
			22: numbervalue = 40'b0000000000111100000000000000000000000000;
			23: numbervalue = 40'b0000000000111100000000000000000000000000;
			24: numbervalue = 40'b0000000000111100000000000000000000000000;
			25: numbervalue = 40'b0000000000111100000000000000000000000000;
			26: numbervalue = 40'b0000000000111100000000000000000000000000;
			27: numbervalue = 40'b0000000000111100000000000000000000000000;
			28: numbervalue = 40'b0000000000111100000000000000000000000000;
			29: numbervalue = 40'b0000000000111111111111111111000000000000;
			30: numbervalue = 40'b0000000000111111111111111111000000000000;
			31: numbervalue = 40'b0000000000111111111111111111000000000000;
			32: numbervalue = 40'b0000000000000000000000000000000000000000;
			33: numbervalue = 40'b0000000000000000000000000000000000000000;
			34: numbervalue = 40'b0000000000000000000000000000000000000000;
			35: numbervalue = 40'b0000000000000000000000000000000000000000;
			36: numbervalue = 40'b0000000000000000000000000000000000000000;
			37: numbervalue = 40'b0000000000000000000000000000000000000000;
			38: numbervalue = 40'b0000000000000000000000000000000000000000;
			39: numbervalue = 40'b0000000000000000000000000000000000000000;
			default: numbervalue = 40'd0;
		endcase 
		
			3'd7:case(row) //1
			0: numbervalue =  40'b0000000000000000000000000000000000000000;
			1: numbervalue =  40'b0000000000000000000000000000000000000000;
			2: numbervalue =  40'b0000000000000000000000000000000000000000;
			3: numbervalue =  40'b0000000000000000000000000000000000000000;
			4: numbervalue =  40'b0000000000000000000000000000000000000000;
			5: numbervalue =  40'b0000000000000000000000000000000000000000;
			6: numbervalue =  40'b0000000000000000000000000000000000000000;
			7: numbervalue =  40'b0000000000000000000000000000000000000000;
			8: numbervalue =  40'b0000000000000000001111000000000000000000;
			9: numbervalue =  40'b0000000000000000011111000000000000000000;
			10: numbervalue=  40'b0000000000000000111111000000000000000000;
			11: numbervalue = 40'b0000000000000001111111000000000000000000;
			12: numbervalue = 40'b0000000000000011111111000000000000000000;
			13: numbervalue = 40'b0000000000000111111111000000000000000000;
			14: numbervalue = 40'b0000000000001110011111000000000000000000;
			15: numbervalue = 40'b0000000000011100011111000000000000000000;
			16: numbervalue = 40'b0000000000000000011111000000000000000000;
			17: numbervalue = 40'b0000000000000000011111000000000000000000;
			18: numbervalue = 40'b0000000000000000011111000000000000000000;
			19: numbervalue = 40'b0000000000000000011111000000000000000000;
			20: numbervalue = 40'b0000000000000000011111000000000000000000;
			21: numbervalue = 40'b0000000000000000011111000000000000000000;
			22: numbervalue = 40'b0000000000000000011111000000000000000000;
			23: numbervalue = 40'b0000000000000000011111000000000000000000;
			24: numbervalue = 40'b0000000000000000011111000000000000000000;
			25: numbervalue = 40'b0000000000000000011111000000000000000000;
			26: numbervalue = 40'b0000000000000000011111000000000000000000;
			27: numbervalue = 40'b0000000000000000011111000000000000000000;
			28: numbervalue = 40'b0000000000000000011111000000000000000000;
			29: numbervalue = 40'b0000000000011111111111111111000000000000;
			30: numbervalue = 40'b0000000000011111111111111111000000000000;
			31: numbervalue = 40'b0000000000011111111111111111000000000000;
			32: numbervalue = 40'b0000000000000000000000000000000000000000;
			33: numbervalue = 40'b0000000000000000000000000000000000000000;
			34: numbervalue = 40'b0000000000000000000000000000000000000000;
			35: numbervalue = 40'b0000000000000000000000000000000000000000;
			36: numbervalue = 40'b0000000000000000000000000000000000000000;
			37: numbervalue = 40'b0000000000000000000000000000000000000000;
			38: numbervalue = 40'b0000000000000000000000000000000000000000;
			39: numbervalue = 40'b0000000000000000000000000000000000000000;
			default: numbervalue = 40'd0;
		endcase
		default: numbervalue = 40'd0;
	endcase
end


endmodule
